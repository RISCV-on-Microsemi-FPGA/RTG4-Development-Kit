`timescale 1ns/10ps
`define RANDOMIZE

module CSRFile(
  input   clk,
  input   reset,
  input   io_prci_reset,
  input   io_prci_id,
  input   io_prci_interrupts_meip,
  input   io_prci_interrupts_seip,
  input   io_prci_interrupts_debug,
  input   io_prci_interrupts_mtip,
  input   io_prci_interrupts_msip,
  input  [11:0] io_rw_addr,
  input  [2:0] io_rw_cmd,
  output [31:0] io_rw_rdata,
  input  [31:0] io_rw_wdata,
  output  io_csr_stall,
  output  io_csr_xcpt,
  output  io_eret,
  output  io_singleStep,
  output  io_status_debug,
  output [1:0] io_status_prv,
  output  io_status_sd,
  output [30:0] io_status_zero3,
  output  io_status_sd_rv32,
  output [1:0] io_status_zero2,
  output [4:0] io_status_vm,
  output [3:0] io_status_zero1,
  output  io_status_mxr,
  output  io_status_pum,
  output  io_status_mprv,
  output [1:0] io_status_xs,
  output [1:0] io_status_fs,
  output [1:0] io_status_mpp,
  output [1:0] io_status_hpp,
  output  io_status_spp,
  output  io_status_mpie,
  output  io_status_hpie,
  output  io_status_spie,
  output  io_status_upie,
  output  io_status_mie,
  output  io_status_hie,
  output  io_status_sie,
  output  io_status_uie,
  output [6:0] io_ptbr_asid,
  output [21:0] io_ptbr_ppn,
  output [31:0] io_evec,
  input   io_exception,
  input   io_retire,
  input  [31:0] io_cause,
  input  [31:0] io_pc,
  input  [31:0] io_badaddr,
  output  io_fatc,
  output [31:0] io_time,
  output [2:0] io_fcsr_rm,
  input   io_fcsr_flags_valid,
  input  [4:0] io_fcsr_flags_bits,
  input   io_rocc_cmd_ready,
  output  io_rocc_cmd_valid,
  output [6:0] io_rocc_cmd_bits_inst_funct,
  output [4:0] io_rocc_cmd_bits_inst_rs2,
  output [4:0] io_rocc_cmd_bits_inst_rs1,
  output  io_rocc_cmd_bits_inst_xd,
  output  io_rocc_cmd_bits_inst_xs1,
  output  io_rocc_cmd_bits_inst_xs2,
  output [4:0] io_rocc_cmd_bits_inst_rd,
  output [6:0] io_rocc_cmd_bits_inst_opcode,
  output [31:0] io_rocc_cmd_bits_rs1,
  output [31:0] io_rocc_cmd_bits_rs2,
  output  io_rocc_cmd_bits_status_debug,
  output [1:0] io_rocc_cmd_bits_status_prv,
  output  io_rocc_cmd_bits_status_sd,
  output [30:0] io_rocc_cmd_bits_status_zero3,
  output  io_rocc_cmd_bits_status_sd_rv32,
  output [1:0] io_rocc_cmd_bits_status_zero2,
  output [4:0] io_rocc_cmd_bits_status_vm,
  output [3:0] io_rocc_cmd_bits_status_zero1,
  output  io_rocc_cmd_bits_status_mxr,
  output  io_rocc_cmd_bits_status_pum,
  output  io_rocc_cmd_bits_status_mprv,
  output [1:0] io_rocc_cmd_bits_status_xs,
  output [1:0] io_rocc_cmd_bits_status_fs,
  output [1:0] io_rocc_cmd_bits_status_mpp,
  output [1:0] io_rocc_cmd_bits_status_hpp,
  output  io_rocc_cmd_bits_status_spp,
  output  io_rocc_cmd_bits_status_mpie,
  output  io_rocc_cmd_bits_status_hpie,
  output  io_rocc_cmd_bits_status_spie,
  output  io_rocc_cmd_bits_status_upie,
  output  io_rocc_cmd_bits_status_mie,
  output  io_rocc_cmd_bits_status_hie,
  output  io_rocc_cmd_bits_status_sie,
  output  io_rocc_cmd_bits_status_uie,
  output  io_rocc_resp_ready,
  input   io_rocc_resp_valid,
  input  [4:0] io_rocc_resp_bits_rd,
  input  [31:0] io_rocc_resp_bits_data,
  output  io_rocc_mem_req_ready,
  input   io_rocc_mem_req_valid,
  input  [31:0] io_rocc_mem_req_bits_addr,
  input  [8:0] io_rocc_mem_req_bits_tag,
  input  [4:0] io_rocc_mem_req_bits_cmd,
  input  [2:0] io_rocc_mem_req_bits_typ,
  input   io_rocc_mem_req_bits_phys,
  input  [31:0] io_rocc_mem_req_bits_data,
  input   io_rocc_mem_s1_kill,
  input  [31:0] io_rocc_mem_s1_data,
  output  io_rocc_mem_s2_nack,
  output  io_rocc_mem_resp_valid,
  output [31:0] io_rocc_mem_resp_bits_addr,
  output [8:0] io_rocc_mem_resp_bits_tag,
  output [4:0] io_rocc_mem_resp_bits_cmd,
  output [2:0] io_rocc_mem_resp_bits_typ,
  output [31:0] io_rocc_mem_resp_bits_data,
  output  io_rocc_mem_resp_bits_replay,
  output  io_rocc_mem_resp_bits_has_data,
  output [31:0] io_rocc_mem_resp_bits_data_word_bypass,
  output [31:0] io_rocc_mem_resp_bits_store_data,
  output  io_rocc_mem_replay_next,
  output  io_rocc_mem_xcpt_ma_ld,
  output  io_rocc_mem_xcpt_ma_st,
  output  io_rocc_mem_xcpt_pf_ld,
  output  io_rocc_mem_xcpt_pf_st,
  input   io_rocc_mem_invalidate_lr,
  output  io_rocc_mem_ordered,
  input   io_rocc_busy,
  input   io_rocc_interrupt,
  output  io_rocc_autl_acquire_ready,
  input   io_rocc_autl_acquire_valid,
  input  [25:0] io_rocc_autl_acquire_bits_addr_block,
  input   io_rocc_autl_acquire_bits_client_xact_id,
  input  [2:0] io_rocc_autl_acquire_bits_addr_beat,
  input   io_rocc_autl_acquire_bits_is_builtin_type,
  input  [2:0] io_rocc_autl_acquire_bits_a_type,
  input  [11:0] io_rocc_autl_acquire_bits_union,
  input  [63:0] io_rocc_autl_acquire_bits_data,
  input   io_rocc_autl_grant_ready,
  output  io_rocc_autl_grant_valid,
  output [2:0] io_rocc_autl_grant_bits_addr_beat,
  output  io_rocc_autl_grant_bits_client_xact_id,
  output [1:0] io_rocc_autl_grant_bits_manager_xact_id,
  output  io_rocc_autl_grant_bits_is_builtin_type,
  output [3:0] io_rocc_autl_grant_bits_g_type,
  output [63:0] io_rocc_autl_grant_bits_data,
  output  io_rocc_fpu_req_ready,
  input   io_rocc_fpu_req_valid,
  input  [4:0] io_rocc_fpu_req_bits_cmd,
  input   io_rocc_fpu_req_bits_ldst,
  input   io_rocc_fpu_req_bits_wen,
  input   io_rocc_fpu_req_bits_ren1,
  input   io_rocc_fpu_req_bits_ren2,
  input   io_rocc_fpu_req_bits_ren3,
  input   io_rocc_fpu_req_bits_swap12,
  input   io_rocc_fpu_req_bits_swap23,
  input   io_rocc_fpu_req_bits_single,
  input   io_rocc_fpu_req_bits_fromint,
  input   io_rocc_fpu_req_bits_toint,
  input   io_rocc_fpu_req_bits_fastpipe,
  input   io_rocc_fpu_req_bits_fma,
  input   io_rocc_fpu_req_bits_div,
  input   io_rocc_fpu_req_bits_sqrt,
  input   io_rocc_fpu_req_bits_round,
  input   io_rocc_fpu_req_bits_wflags,
  input  [2:0] io_rocc_fpu_req_bits_rm,
  input  [1:0] io_rocc_fpu_req_bits_typ,
  input  [64:0] io_rocc_fpu_req_bits_in1,
  input  [64:0] io_rocc_fpu_req_bits_in2,
  input  [64:0] io_rocc_fpu_req_bits_in3,
  input   io_rocc_fpu_resp_ready,
  output  io_rocc_fpu_resp_valid,
  output [64:0] io_rocc_fpu_resp_bits_data,
  output [4:0] io_rocc_fpu_resp_bits_exc,
  output  io_rocc_exception,
  output [11:0] io_rocc_csr_waddr,
  output [31:0] io_rocc_csr_wdata,
  output  io_rocc_csr_wen,
  output  io_rocc_host_id,
  output  io_interrupt,
  output [31:0] io_interrupt_cause,
  output [3:0] io_bp_0_control_tdrtype,
  output [4:0] io_bp_0_control_bpamaskmax,
  output [3:0] io_bp_0_control_reserved,
  output [7:0] io_bp_0_control_bpaction,
  output [3:0] io_bp_0_control_bpmatch,
  output  io_bp_0_control_m,
  output  io_bp_0_control_h,
  output  io_bp_0_control_s,
  output  io_bp_0_control_u,
  output  io_bp_0_control_r,
  output  io_bp_0_control_w,
  output  io_bp_0_control_x,
  output [31:0] io_bp_0_address,
  output [3:0] io_bp_1_control_tdrtype,
  output [4:0] io_bp_1_control_bpamaskmax,
  output [3:0] io_bp_1_control_reserved,
  output [7:0] io_bp_1_control_bpaction,
  output [3:0] io_bp_1_control_bpmatch,
  output  io_bp_1_control_m,
  output  io_bp_1_control_h,
  output  io_bp_1_control_s,
  output  io_bp_1_control_u,
  output  io_bp_1_control_r,
  output  io_bp_1_control_w,
  output  io_bp_1_control_x,
  output [31:0] io_bp_1_address
);
  wire  T_5012_debug;
  wire [1:0] T_5012_prv;
  wire  T_5012_sd;
  wire [30:0] T_5012_zero3;
  wire  T_5012_sd_rv32;
  wire [1:0] T_5012_zero2;
  wire [4:0] T_5012_vm;
  wire [3:0] T_5012_zero1;
  wire  T_5012_mxr;
  wire  T_5012_pum;
  wire  T_5012_mprv;
  wire [1:0] T_5012_xs;
  wire [1:0] T_5012_fs;
  wire [1:0] T_5012_mpp;
  wire [1:0] T_5012_hpp;
  wire  T_5012_spp;
  wire  T_5012_mpie;
  wire  T_5012_hpie;
  wire  T_5012_spie;
  wire  T_5012_upie;
  wire  T_5012_mie;
  wire  T_5012_hie;
  wire  T_5012_sie;
  wire  T_5012_uie;
  wire [66:0] T_5038;
  wire  T_5039;
  wire  T_5040;
  wire  T_5041;
  wire  T_5042;
  wire  T_5043;
  wire  T_5044;
  wire  T_5045;
  wire  T_5046;
  wire  T_5047;
  wire [1:0] T_5048;
  wire [1:0] T_5049;
  wire [1:0] T_5050;
  wire [1:0] T_5051;
  wire  T_5052;
  wire  T_5053;
  wire  T_5054;
  wire [3:0] T_5055;
  wire [4:0] T_5056;
  wire [1:0] T_5057;
  wire  T_5058;
  wire [30:0] T_5059;
  wire  T_5060;
  wire [1:0] T_5061;
  wire  T_5062;
  wire  reset_mstatus_debug;
  wire [1:0] reset_mstatus_prv;
  wire  reset_mstatus_sd;
  wire [30:0] reset_mstatus_zero3;
  wire  reset_mstatus_sd_rv32;
  wire [1:0] reset_mstatus_zero2;
  wire [4:0] reset_mstatus_vm;
  wire [3:0] reset_mstatus_zero1;
  wire  reset_mstatus_mxr;
  wire  reset_mstatus_pum;
  wire  reset_mstatus_mprv;
  wire [1:0] reset_mstatus_xs;
  wire [1:0] reset_mstatus_fs;
  wire [1:0] reset_mstatus_mpp;
  wire [1:0] reset_mstatus_hpp;
  wire  reset_mstatus_spp;
  wire  reset_mstatus_mpie;
  wire  reset_mstatus_hpie;
  wire  reset_mstatus_spie;
  wire  reset_mstatus_upie;
  wire  reset_mstatus_mie;
  wire  reset_mstatus_hie;
  wire  reset_mstatus_sie;
  wire  reset_mstatus_uie;
  reg  reg_mstatus_debug;
  reg [31:0] GEN_152;
  reg [1:0] reg_mstatus_prv;
  reg [31:0] GEN_153;
  reg  reg_mstatus_sd;
  reg [31:0] GEN_154;
  reg [30:0] reg_mstatus_zero3;
  reg [31:0] GEN_155;
  reg  reg_mstatus_sd_rv32;
  reg [31:0] GEN_156;
  reg [1:0] reg_mstatus_zero2;
  reg [31:0] GEN_157;
  reg [4:0] reg_mstatus_vm;
  reg [31:0] GEN_158;
  reg [3:0] reg_mstatus_zero1;
  reg [31:0] GEN_159;
  reg  reg_mstatus_mxr;
  reg [31:0] GEN_160;
  reg  reg_mstatus_pum;
  reg [31:0] GEN_161;
  reg  reg_mstatus_mprv;
  reg [31:0] GEN_162;
  reg [1:0] reg_mstatus_xs;
  reg [31:0] GEN_163;
  reg [1:0] reg_mstatus_fs;
  reg [31:0] GEN_164;
  reg [1:0] reg_mstatus_mpp;
  reg [31:0] GEN_165;
  reg [1:0] reg_mstatus_hpp;
  reg [31:0] GEN_166;
  reg  reg_mstatus_spp;
  reg [31:0] GEN_167;
  reg  reg_mstatus_mpie;
  reg [31:0] GEN_168;
  reg  reg_mstatus_hpie;
  reg [31:0] GEN_175;
  reg  reg_mstatus_spie;
  reg [31:0] GEN_176;
  reg  reg_mstatus_upie;
  reg [31:0] GEN_177;
  reg  reg_mstatus_mie;
  reg [31:0] GEN_178;
  reg  reg_mstatus_hie;
  reg [31:0] GEN_179;
  reg  reg_mstatus_sie;
  reg [31:0] GEN_180;
  reg  reg_mstatus_uie;
  reg [31:0] GEN_181;
  wire [1:0] T_5150_xdebugver;
  wire  T_5150_ndreset;
  wire  T_5150_fullreset;
  wire [11:0] T_5150_hwbpcount;
  wire  T_5150_ebreakm;
  wire  T_5150_ebreakh;
  wire  T_5150_ebreaks;
  wire  T_5150_ebreaku;
  wire  T_5150_zero2;
  wire  T_5150_stopcycle;
  wire  T_5150_stoptime;
  wire [2:0] T_5150_cause;
  wire  T_5150_debugint;
  wire  T_5150_zero1;
  wire  T_5150_halt;
  wire  T_5150_step;
  wire [1:0] T_5150_prv;
  wire [31:0] T_5169;
  wire [1:0] T_5170;
  wire  T_5171;
  wire  T_5172;
  wire  T_5173;
  wire  T_5174;
  wire [2:0] T_5175;
  wire  T_5176;
  wire  T_5177;
  wire  T_5178;
  wire  T_5179;
  wire  T_5180;
  wire  T_5181;
  wire  T_5182;
  wire [11:0] T_5183;
  wire  T_5184;
  wire  T_5185;
  wire [1:0] T_5186;
  wire [1:0] reset_dcsr_xdebugver;
  wire  reset_dcsr_ndreset;
  wire  reset_dcsr_fullreset;
  wire [11:0] reset_dcsr_hwbpcount;
  wire  reset_dcsr_ebreakm;
  wire  reset_dcsr_ebreakh;
  wire  reset_dcsr_ebreaks;
  wire  reset_dcsr_ebreaku;
  wire  reset_dcsr_zero2;
  wire  reset_dcsr_stopcycle;
  wire  reset_dcsr_stoptime;
  wire [2:0] reset_dcsr_cause;
  wire  reset_dcsr_debugint;
  wire  reset_dcsr_zero1;
  wire  reset_dcsr_halt;
  wire  reset_dcsr_step;
  wire [1:0] reset_dcsr_prv;
  reg [1:0] reg_dcsr_xdebugver;
  reg [31:0] GEN_182;
  reg  reg_dcsr_ndreset;
  reg [31:0] GEN_185;
  reg  reg_dcsr_fullreset;
  reg [31:0] GEN_186;
  reg [11:0] reg_dcsr_hwbpcount;
  reg [31:0] GEN_187;
  reg  reg_dcsr_ebreakm;
  reg [31:0] GEN_188;
  reg  reg_dcsr_ebreakh;
  reg [31:0] GEN_189;
  reg  reg_dcsr_ebreaks;
  reg [31:0] GEN_190;
  reg  reg_dcsr_ebreaku;
  reg [31:0] GEN_191;
  reg  reg_dcsr_zero2;
  reg [31:0] GEN_192;
  reg  reg_dcsr_stopcycle;
  reg [31:0] GEN_201;
  reg  reg_dcsr_stoptime;
  reg [31:0] GEN_202;
  reg [2:0] reg_dcsr_cause;
  reg [31:0] GEN_203;
  reg  reg_dcsr_debugint;
  reg [31:0] GEN_204;
  reg  reg_dcsr_zero1;
  reg [31:0] GEN_205;
  reg  reg_dcsr_halt;
  reg [31:0] GEN_206;
  reg  reg_dcsr_step;
  reg [31:0] GEN_207;
  reg [1:0] reg_dcsr_prv;
  reg [31:0] GEN_208;
  wire  T_5252_rocc;
  wire  T_5252_meip;
  wire  T_5252_heip;
  wire  T_5252_seip;
  wire  T_5252_ueip;
  wire  T_5252_mtip;
  wire  T_5252_htip;
  wire  T_5252_stip;
  wire  T_5252_utip;
  wire  T_5252_msip;
  wire  T_5252_hsip;
  wire  T_5252_ssip;
  wire  T_5252_usip;
  wire [12:0] T_5267;
  wire  T_5268;
  wire  T_5269;
  wire  T_5270;
  wire  T_5271;
  wire  T_5272;
  wire  T_5273;
  wire  T_5274;
  wire  T_5275;
  wire  T_5276;
  wire  T_5277;
  wire  T_5278;
  wire  T_5279;
  wire  T_5280;
  wire  T_5281_rocc;
  wire  T_5281_meip;
  wire  T_5281_heip;
  wire  T_5281_seip;
  wire  T_5281_ueip;
  wire  T_5281_mtip;
  wire  T_5281_htip;
  wire  T_5281_stip;
  wire  T_5281_utip;
  wire  T_5281_msip;
  wire  T_5281_hsip;
  wire  T_5281_ssip;
  wire  T_5281_usip;
  wire  T_5302_rocc;
  wire  T_5302_meip;
  wire  T_5302_heip;
  wire  T_5302_seip;
  wire  T_5302_ueip;
  wire  T_5302_mtip;
  wire  T_5302_htip;
  wire  T_5302_stip;
  wire  T_5302_utip;
  wire  T_5302_msip;
  wire  T_5302_hsip;
  wire  T_5302_ssip;
  wire  T_5302_usip;
  wire [1:0] T_5319;
  wire [2:0] T_5320;
  wire [1:0] T_5321;
  wire [2:0] T_5322;
  wire [5:0] T_5323;
  wire [1:0] T_5324;
  wire [2:0] T_5325;
  wire [1:0] T_5326;
  wire [1:0] T_5327;
  wire [3:0] T_5328;
  wire [6:0] T_5329;
  wire [12:0] supported_interrupts;
  wire  exception;
  reg  reg_debug;
  reg [31:0] GEN_209;
  reg [31:0] reg_dpc;
  reg [31:0] GEN_210;
  reg [31:0] reg_dscratch;
  reg [31:0] GEN_211;
  reg  reg_singleStepped;
  reg [31:0] GEN_212;
  wire  T_5346;
  wire  GEN_27;
  wire  T_5349;
  wire  GEN_28;
  wire  T_5360;
  wire  T_5362;
  wire  T_5363;
  wire  T_5364;
  wire  T_5366;
  reg  reg_tdrselect_tdrmode;
  reg [31:0] GEN_213;
  reg [29:0] reg_tdrselect_reserved;
  reg [31:0] GEN_214;
  reg  reg_tdrselect_tdrindex;
  reg [31:0] GEN_215;
  reg [3:0] reg_bp_0_control_tdrtype;
  reg [31:0] GEN_216;
  reg [4:0] reg_bp_0_control_bpamaskmax;
  reg [31:0] GEN_217;
  reg [3:0] reg_bp_0_control_reserved;
  reg [31:0] GEN_218;
  reg [7:0] reg_bp_0_control_bpaction;
  reg [31:0] GEN_219;
  reg [3:0] reg_bp_0_control_bpmatch;
  reg [31:0] GEN_220;
  reg  reg_bp_0_control_m;
  reg [31:0] GEN_221;
  reg  reg_bp_0_control_h;
  reg [31:0] GEN_222;
  reg  reg_bp_0_control_s;
  reg [31:0] GEN_223;
  reg  reg_bp_0_control_u;
  reg [31:0] GEN_224;
  reg  reg_bp_0_control_r;
  reg [31:0] GEN_225;
  reg  reg_bp_0_control_w;
  reg [31:0] GEN_228;
  reg  reg_bp_0_control_x;
  reg [31:0] GEN_229;
  reg [31:0] reg_bp_0_address;
  reg [31:0] GEN_230;
  reg [3:0] reg_bp_1_control_tdrtype;
  reg [31:0] GEN_231;
  reg [4:0] reg_bp_1_control_bpamaskmax;
  reg [31:0] GEN_232;
  reg [3:0] reg_bp_1_control_reserved;
  reg [31:0] GEN_233;
  reg [7:0] reg_bp_1_control_bpaction;
  reg [31:0] GEN_234;
  reg [3:0] reg_bp_1_control_bpmatch;
  reg [31:0] GEN_235;
  reg  reg_bp_1_control_m;
  reg [31:0] GEN_236;
  reg  reg_bp_1_control_h;
  reg [31:0] GEN_237;
  reg  reg_bp_1_control_s;
  reg [31:0] GEN_238;
  reg  reg_bp_1_control_u;
  reg [31:0] GEN_239;
  reg  reg_bp_1_control_r;
  reg [31:0] GEN_240;
  reg  reg_bp_1_control_w;
  reg [31:0] GEN_243;
  reg  reg_bp_1_control_x;
  reg [31:0] GEN_246;
  reg [31:0] reg_bp_1_address;
  reg [31:0] GEN_249;
  reg [31:0] reg_mie;
  reg [31:0] GEN_252;
  reg [31:0] reg_mideleg;
  reg [31:0] GEN_255;
  reg [31:0] reg_medeleg;
  reg [31:0] GEN_256;
  reg  reg_mip_rocc;
  reg [31:0] GEN_257;
  reg  reg_mip_meip;
  reg [31:0] GEN_258;
  reg  reg_mip_heip;
  reg [31:0] GEN_259;
  reg  reg_mip_seip;
  reg [31:0] GEN_260;
  reg  reg_mip_ueip;
  reg [31:0] GEN_261;
  reg  reg_mip_mtip;
  reg [31:0] GEN_262;
  reg  reg_mip_htip;
  reg [31:0] GEN_263;
  reg  reg_mip_stip;
  reg [31:0] GEN_264;
  reg  reg_mip_utip;
  reg [31:0] GEN_265;
  reg  reg_mip_msip;
  reg [31:0] GEN_266;
  reg  reg_mip_hsip;
  reg [31:0] GEN_267;
  reg  reg_mip_ssip;
  reg [31:0] GEN_268;
  reg  reg_mip_usip;
  reg [31:0] GEN_269;
  reg [31:0] reg_mepc;
  reg [31:0] GEN_270;
  reg [31:0] reg_mcause;
  reg [31:0] GEN_271;
  reg [31:0] reg_mbadaddr;
  reg [31:0] GEN_272;
  reg [31:0] reg_mscratch;
  reg [31:0] GEN_273;
  reg [31:0] reg_mtvec;
  reg [31:0] GEN_274;
  reg [31:0] reg_sepc;
  reg [31:0] GEN_275;
  reg [31:0] reg_scause;
  reg [31:0] GEN_276;
  reg [31:0] reg_sbadaddr;
  reg [31:0] GEN_277;
  reg [31:0] reg_sscratch;
  reg [31:0] GEN_278;
  reg [31:0] reg_stvec;
  reg [31:0] GEN_279;
  reg [6:0] reg_sptbr_asid;
  reg [31:0] GEN_282;
  reg [21:0] reg_sptbr_ppn;
  reg [31:0] GEN_283;
  reg  reg_wfi;
  reg [31:0] GEN_284;
  reg [4:0] reg_fflags;
  reg [31:0] GEN_285;
  reg [2:0] reg_frm;
  reg [31:0] GEN_286;
  reg [5:0] T_5570;
  reg [31:0] GEN_287;
  wire [5:0] GEN_437;
  wire [6:0] T_5571;
  reg [57:0] T_5573;
  reg [63:0] GEN_288;
  wire  T_5574;
  wire [58:0] T_5576;
  wire [57:0] T_5577;
  wire [57:0] GEN_29;
  wire [63:0] T_5578;
  reg [5:0] T_5581;
  reg [31:0] GEN_289;
  wire [6:0] T_5582;
  reg [57:0] T_5584;
  reg [63:0] GEN_290;
  wire  T_5585;
  wire [58:0] T_5587;
  wire [57:0] T_5588;
  wire [57:0] GEN_30;
  wire [63:0] reg_cycle;
  wire  mip_rocc;
  wire  mip_meip;
  wire  mip_heip;
  wire  mip_seip;
  wire  mip_ueip;
  wire  mip_mtip;
  wire  mip_htip;
  wire  mip_stip;
  wire  mip_utip;
  wire  mip_msip;
  wire  mip_hsip;
  wire  mip_ssip;
  wire  mip_usip;
  wire [1:0] T_5602;
  wire [2:0] T_5603;
  wire [1:0] T_5604;
  wire [2:0] T_5605;
  wire [5:0] T_5606;
  wire [1:0] T_5607;
  wire [2:0] T_5608;
  wire [1:0] T_5609;
  wire [1:0] T_5610;
  wire [3:0] T_5611;
  wire [6:0] T_5612;
  wire [12:0] T_5613;
  wire [12:0] read_mip;
  wire [31:0] GEN_438;
  wire [31:0] pending_interrupts;
  wire  T_5615;
  wire  T_5617;
  wire  T_5619;
  wire  T_5620;
  wire  T_5621;
  wire  T_5622;
  wire [31:0] T_5623;
  wire [31:0] T_5624;
  wire [31:0] m_interrupts;
  wire  T_5629;
  wire  T_5631;
  wire  T_5632;
  wire  T_5633;
  wire  T_5634;
  wire [31:0] T_5635;
  wire [31:0] s_interrupts;
  wire [31:0] all_interrupts;
  wire  T_5638;
  wire  T_5639;
  wire  T_5640;
  wire  T_5641;
  wire  T_5642;
  wire  T_5643;
  wire  T_5644;
  wire  T_5645;
  wire  T_5646;
  wire  T_5647;
  wire  T_5648;
  wire  T_5649;
  wire  T_5650;
  wire  T_5651;
  wire  T_5652;
  wire  T_5653;
  wire  T_5654;
  wire  T_5655;
  wire  T_5656;
  wire  T_5657;
  wire  T_5658;
  wire  T_5659;
  wire  T_5660;
  wire  T_5661;
  wire  T_5662;
  wire  T_5663;
  wire  T_5664;
  wire  T_5665;
  wire  T_5666;
  wire  T_5667;
  wire  T_5668;
  wire [4:0] T_5702;
  wire [4:0] T_5703;
  wire [4:0] T_5704;
  wire [4:0] T_5705;
  wire [4:0] T_5706;
  wire [4:0] T_5707;
  wire [4:0] T_5708;
  wire [4:0] T_5709;
  wire [4:0] T_5710;
  wire [4:0] T_5711;
  wire [4:0] T_5712;
  wire [4:0] T_5713;
  wire [4:0] T_5714;
  wire [4:0] T_5715;
  wire [4:0] T_5716;
  wire [4:0] T_5717;
  wire [4:0] T_5718;
  wire [4:0] T_5719;
  wire [4:0] T_5720;
  wire [4:0] T_5721;
  wire [4:0] T_5722;
  wire [4:0] T_5723;
  wire [4:0] T_5724;
  wire [4:0] T_5725;
  wire [4:0] T_5726;
  wire [4:0] T_5727;
  wire [4:0] T_5728;
  wire [4:0] T_5729;
  wire [4:0] T_5730;
  wire [4:0] T_5731;
  wire [4:0] T_5732;
  wire [31:0] GEN_439;
  wire [32:0] T_5733;
  wire [31:0] interruptCause;
  wire  T_5735;
  wire  T_5738;
  wire  T_5739;
  wire  T_5744;
  wire  GEN_31;
  wire [31:0] GEN_32;
  wire  system_insn;
  wire  T_5747;
  wire  T_5749;
  wire  cpu_ren;
  wire [1:0] T_5750;
  wire [2:0] T_5751;
  wire [1:0] T_5752;
  wire [2:0] T_5753;
  wire [5:0] T_5754;
  wire [1:0] T_5755;
  wire [2:0] T_5756;
  wire [3:0] T_5757;
  wire [5:0] T_5758;
  wire [8:0] T_5759;
  wire [14:0] T_5760;
  wire [1:0] T_5761;
  wire [3:0] T_5762;
  wire [8:0] T_5763;
  wire [9:0] T_5764;
  wire [13:0] T_5765;
  wire [31:0] T_5766;
  wire [33:0] T_5767;
  wire [2:0] T_5768;
  wire [3:0] T_5769;
  wire [37:0] T_5770;
  wire [51:0] T_5771;
  wire [66:0] T_5772;
  wire [31:0] read_mstatus;
  wire [30:0] T_5773;
  wire [31:0] T_5774;
  wire  GEN_0;
  wire  GEN_33;
  wire  GEN_1;
  wire  GEN_34;
  wire [1:0] T_5789;
  wire  GEN_2;
  wire  GEN_35;
  wire [2:0] T_5790;
  wire  GEN_3;
  wire  GEN_36;
  wire  GEN_4;
  wire  GEN_37;
  wire [1:0] T_5791;
  wire  GEN_5;
  wire  GEN_38;
  wire [2:0] T_5792;
  wire [5:0] T_5793;
  wire [7:0] GEN_6;
  wire [7:0] GEN_39;
  wire [3:0] GEN_7;
  wire [3:0] GEN_40;
  wire [11:0] T_5794;
  wire  GEN_8;
  wire  GEN_41;
  wire [12:0] T_5795;
  wire [3:0] GEN_9;
  wire [3:0] GEN_42;
  wire [4:0] GEN_10;
  wire [4:0] GEN_43;
  wire [8:0] T_5796;
  wire [3:0] GEN_11;
  wire [3:0] GEN_44;
  wire [12:0] T_5797;
  wire [25:0] T_5798;
  wire [31:0] T_5799;
  wire [2:0] T_5822;
  wire [1:0] T_5823;
  wire [4:0] T_5824;
  wire [3:0] T_5825;
  wire [1:0] T_5826;
  wire [5:0] T_5827;
  wire [10:0] T_5828;
  wire [1:0] T_5829;
  wire [1:0] T_5830;
  wire [3:0] T_5831;
  wire [12:0] T_5832;
  wire [2:0] T_5833;
  wire [3:0] T_5834;
  wire [16:0] T_5835;
  wire [20:0] T_5836;
  wire [31:0] T_5837;
  wire [31:0] T_5838;
  wire [31:0] T_5839;
  wire  T_5844;
  wire  T_5846;
  wire  T_5848;
  wire  T_5850;
  wire  T_5852;
  wire  T_5854;
  wire  T_5856;
  wire  T_5858;
  wire  T_5860;
  wire  T_5862;
  wire  T_5864;
  wire  T_5866;
  wire  T_5868;
  wire  T_5870;
  wire  T_5872;
  wire  T_5874;
  wire  T_5876;
  wire  T_5878;
  wire  T_5880;
  wire  T_5882;
  wire  T_5884;
  wire  T_5886;
  wire  T_5888;
  wire  T_5890;
  wire  T_5892;
  wire  T_5894;
  wire  T_5896;
  wire  T_5898;
  wire  T_5900;
  wire  T_5902;
  wire  T_5904;
  wire  T_5906;
  wire  T_5907;
  wire  T_5908;
  wire  T_5909;
  wire  T_5910;
  wire  T_5911;
  wire  T_5912;
  wire  T_5913;
  wire  T_5914;
  wire  T_5915;
  wire  T_5916;
  wire  T_5917;
  wire  T_5918;
  wire  T_5919;
  wire  T_5920;
  wire  T_5921;
  wire  T_5922;
  wire  T_5923;
  wire  T_5924;
  wire  T_5925;
  wire  T_5926;
  wire  T_5927;
  wire  T_5928;
  wire  T_5929;
  wire  T_5930;
  wire  T_5931;
  wire  T_5932;
  wire  T_5933;
  wire  T_5934;
  wire  T_5935;
  wire  T_5936;
  wire  addr_valid;
  wire  T_5938;
  wire [1:0] T_5939;
  wire [1:0] T_5940;
  wire  T_5942;
  wire [1:0] T_5943;
  wire [2:0] csr_addr_priv;
  wire [2:0] T_5944;
  wire  priv_sufficient;
  wire [1:0] T_5945;
  wire [1:0] T_5946;
  wire  read_only;
  wire  T_5948;
  wire  T_5949;
  wire  cpu_wen;
  wire  T_5951;
  wire  wen;
  wire  T_5952;
  wire  T_5953;
  wire  T_5954;
  wire [31:0] T_5956;
  wire  T_5957;
  wire [31:0] T_5959;
  wire [31:0] T_5960;
  wire [31:0] T_5963;
  wire [31:0] T_5964;
  wire [31:0] wdata;
  wire  do_system_insn;
  wire [2:0] T_5966;
  wire [7:0] opcode;
  wire  T_5967;
  wire  insn_call;
  wire  T_5968;
  wire  insn_break;
  wire  T_5969;
  wire  insn_ret;
  wire  T_5970;
  wire  insn_sfence_vm;
  wire  T_5971;
  wire  insn_wfi;
  wire  T_5972;
  wire  T_5974;
  wire  T_5976;
  wire  T_5977;
  wire  T_5984;
  wire  T_5985;
  wire  T_5988;
  wire  T_5989;
  wire  T_5990;
  wire  T_5991;
  wire  GEN_45;
  wire  T_5994;
  wire  GEN_46;
  wire  T_5997;
  wire [3:0] GEN_440;
  wire [4:0] T_5999;
  wire [3:0] T_6000;
  wire [1:0] T_6003;
  wire [3:0] T_6004;
  wire [31:0] cause;
  wire [4:0] cause_lsbs;
  wire  T_6005;
  wire  T_6007;
  wire  causeIsDebugInt;
  wire  T_6009;
  wire [1:0] T_6010;
  wire [1:0] T_6011;
  wire [3:0] T_6012;
  wire [3:0] T_6013;
  wire  T_6014;
  wire  causeIsDebugBreak;
  wire  T_6016;
  wire  T_6017;
  wire  T_6018;
  wire [11:0] debugTVec;
  wire [31:0] tvec;
  wire [31:0] epc;
  wire [31:0] T_6038;
  wire  T_6041;
  wire [1:0] T_6042;
  wire  T_6044;
  wire [1:0] T_6045;
  wire  T_6047;
  wire  T_6048;
  wire [31:0] T_6049;
  wire [31:0] T_6051;
  wire [31:0] T_6052;
  wire [31:0] T_6053;
  wire  T_6054;
  wire [1:0] T_6059;
  wire [2:0] T_6060;
  wire  GEN_47;
  wire [31:0] GEN_48;
  wire [2:0] GEN_49;
  wire [1:0] GEN_50;
  wire  T_6062;
  wire [1:0] GEN_55;
  wire [31:0] GEN_58;
  wire [31:0] GEN_59;
  wire [31:0] GEN_60;
  wire  GEN_61;
  wire  GEN_63;
  wire  GEN_65;
  wire [31:0] GEN_66;
  wire [2:0] GEN_67;
  wire [1:0] GEN_68;
  wire [1:0] GEN_73;
  wire [31:0] GEN_76;
  wire [31:0] GEN_77;
  wire [31:0] GEN_78;
  wire  GEN_79;
  wire  GEN_81;
  wire  GEN_88;
  wire  T_6088;
  wire  T_6090;
  wire  GEN_89;
  wire  GEN_91;
  wire  GEN_93;
  wire  GEN_100;
  wire  GEN_101;
  wire  GEN_102;
  wire [1:0] T_6101;
  wire [1:0] GEN_441;
  wire [2:0] T_6102;
  wire [1:0] T_6103;
  wire [2:0] T_6104;
  wire [2:0] GEN_442;
  wire [3:0] T_6105;
  wire [2:0] T_6106;
  wire  T_6108;
  wire  T_6109;
  wire  T_6111;
  wire [31:0] T_6113;
  wire [31:0] T_6115;
  wire [31:0] GEN_12;
  wire [31:0] GEN_104;
  wire [31:0] T_6117;
  wire [63:0] T_6125;
  wire [63:0] T_6127;
  wire [30:0] T_6137;
  wire [31:0] T_6139;
  wire [31:0] T_6141;
  wire [12:0] T_6143;
  wire [31:0] T_6145;
  wire [31:0] T_6147;
  wire [31:0] T_6149;
  wire [31:0] T_6151;
  wire [31:0] T_6153;
  wire [31:0] T_6155;
  wire [31:0] T_6157;
  wire  T_6159;
  wire [31:0] T_6161;
  wire [31:0] T_6163;
  wire [31:0] T_6165;
  wire [31:0] T_6167;
  wire [31:0] T_6169;
  wire [31:0] T_6177;
  wire [31:0] T_6178;
  wire [63:0] GEN_443;
  wire [63:0] T_6182;
  wire [63:0] T_6183;
  wire [63:0] GEN_444;
  wire [63:0] T_6188;
  wire [63:0] GEN_445;
  wire [63:0] T_6189;
  wire [63:0] GEN_446;
  wire [63:0] T_6190;
  wire [63:0] GEN_447;
  wire [63:0] T_6191;
  wire [63:0] GEN_448;
  wire [63:0] T_6192;
  wire [63:0] GEN_449;
  wire [63:0] T_6193;
  wire [63:0] GEN_450;
  wire [63:0] T_6194;
  wire [63:0] GEN_451;
  wire [63:0] T_6195;
  wire [63:0] GEN_452;
  wire [63:0] T_6196;
  wire [63:0] GEN_453;
  wire [63:0] T_6197;
  wire [63:0] GEN_454;
  wire [63:0] T_6198;
  wire [63:0] GEN_455;
  wire [63:0] T_6199;
  wire [63:0] GEN_456;
  wire [63:0] T_6200;
  wire [63:0] GEN_457;
  wire [63:0] T_6201;
  wire [63:0] GEN_458;
  wire [63:0] T_6202;
  wire [63:0] GEN_459;
  wire [63:0] T_6203;
  wire [63:0] GEN_460;
  wire [63:0] T_6204;
  wire [63:0] T_6208;
  wire [4:0] T_6209;
  wire [4:0] GEN_105;
  wire [1:0] supportedModes_0;
  wire  T_6267_debug;
  wire [1:0] T_6267_prv;
  wire  T_6267_sd;
  wire [30:0] T_6267_zero3;
  wire  T_6267_sd_rv32;
  wire [1:0] T_6267_zero2;
  wire [4:0] T_6267_vm;
  wire [3:0] T_6267_zero1;
  wire  T_6267_mxr;
  wire  T_6267_pum;
  wire  T_6267_mprv;
  wire [1:0] T_6267_xs;
  wire [1:0] T_6267_fs;
  wire [1:0] T_6267_mpp;
  wire [1:0] T_6267_hpp;
  wire  T_6267_spp;
  wire  T_6267_mpie;
  wire  T_6267_hpie;
  wire  T_6267_spie;
  wire  T_6267_upie;
  wire  T_6267_mie;
  wire  T_6267_hie;
  wire  T_6267_sie;
  wire  T_6267_uie;
  wire [66:0] T_6293;
  wire  T_6294;
  wire  T_6295;
  wire  T_6296;
  wire  T_6297;
  wire  T_6298;
  wire  T_6299;
  wire  T_6300;
  wire  T_6301;
  wire  T_6302;
  wire [1:0] T_6303;
  wire [1:0] T_6304;
  wire [1:0] T_6305;
  wire [1:0] T_6306;
  wire  T_6307;
  wire  T_6308;
  wire  T_6309;
  wire [3:0] T_6310;
  wire [4:0] T_6311;
  wire [1:0] T_6312;
  wire  T_6313;
  wire [30:0] T_6314;
  wire  T_6315;
  wire [1:0] T_6316;
  wire  T_6317;
  wire  GEN_131;
  wire  GEN_132;
  wire  T_6346_rocc;
  wire  T_6346_meip;
  wire  T_6346_heip;
  wire  T_6346_seip;
  wire  T_6346_ueip;
  wire  T_6346_mtip;
  wire  T_6346_htip;
  wire  T_6346_stip;
  wire  T_6346_utip;
  wire  T_6346_msip;
  wire  T_6346_hsip;
  wire  T_6346_ssip;
  wire  T_6346_usip;
  wire  T_6360;
  wire  T_6361;
  wire  T_6362;
  wire  T_6363;
  wire  T_6364;
  wire  T_6365;
  wire  T_6366;
  wire  T_6367;
  wire  T_6368;
  wire  T_6369;
  wire  T_6370;
  wire  T_6371;
  wire  T_6372;
  wire [31:0] GEN_461;
  wire [31:0] T_6373;
  wire [31:0] GEN_146;
  wire [31:0] T_6374;
  wire [31:0] T_6376;
  wire [31:0] T_6377;
  wire [31:0] GEN_147;
  wire [31:0] GEN_148;
  wire [29:0] T_6378;
  wire [31:0] GEN_462;
  wire [31:0] T_6379;
  wire [31:0] GEN_149;
  wire [31:0] T_6381;
  wire [31:0] GEN_150;
  wire [31:0] GEN_151;
  wire [1:0] T_6419_xdebugver;
  wire  T_6419_ndreset;
  wire  T_6419_fullreset;
  wire [11:0] T_6419_hwbpcount;
  wire  T_6419_ebreakm;
  wire  T_6419_ebreakh;
  wire  T_6419_ebreaks;
  wire  T_6419_ebreaku;
  wire  T_6419_zero2;
  wire  T_6419_stopcycle;
  wire  T_6419_stoptime;
  wire [2:0] T_6419_cause;
  wire  T_6419_debugint;
  wire  T_6419_zero1;
  wire  T_6419_halt;
  wire  T_6419_step;
  wire [1:0] T_6419_prv;
  wire [1:0] T_6437;
  wire [2:0] T_6442;
  wire  T_6447;
  wire  T_6448;
  wire  T_6449;
  wire [11:0] T_6450;
  wire  T_6451;
  wire  T_6452;
  wire [1:0] T_6453;
  wire  GEN_169;
  wire  GEN_170;
  wire  GEN_171;
  wire [31:0] GEN_172;
  wire [31:0] GEN_173;
  wire  T_6466_tdrmode;
  wire [29:0] T_6466_reserved;
  wire  T_6466_tdrindex;
  wire [29:0] T_6471;
  wire  T_6472;
  wire  GEN_174;
  wire  T_6473;
  wire [3:0] T_6500_tdrtype;
  wire [4:0] T_6500_bpamaskmax;
  wire [3:0] T_6500_reserved;
  wire [7:0] T_6500_bpaction;
  wire [3:0] T_6500_bpmatch;
  wire  T_6500_m;
  wire  T_6500_h;
  wire  T_6500_s;
  wire  T_6500_u;
  wire  T_6500_r;
  wire  T_6500_w;
  wire  T_6500_x;
  wire [3:0] T_6520;
  wire [7:0] T_6521;
  wire [3:0] T_6522;
  wire [4:0] T_6523;
  wire [3:0] T_6524;
  wire [3:0] GEN_13;
  wire [4:0] GEN_14;
  wire [3:0] GEN_15;
  wire [7:0] GEN_16;
  wire [3:0] GEN_17;
  wire [3:0] GEN_183;
  wire [3:0] GEN_184;
  wire  GEN_18;
  wire  GEN_19;
  wire  GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire  GEN_193;
  wire  GEN_194;
  wire  GEN_23;
  wire  GEN_195;
  wire  GEN_196;
  wire  GEN_24;
  wire  GEN_197;
  wire  GEN_198;
  wire [3:0] T_6554;
  wire [3:0] GEN_25;
  wire [3:0] GEN_199;
  wire [3:0] GEN_200;
  wire [3:0] GEN_226;
  wire [3:0] GEN_227;
  wire  GEN_241;
  wire  GEN_242;
  wire  GEN_244;
  wire  GEN_245;
  wire  GEN_247;
  wire  GEN_248;
  wire [31:0] GEN_26;
  wire [31:0] GEN_250;
  wire [31:0] GEN_251;
  wire [31:0] GEN_253;
  wire [31:0] GEN_254;
  wire [3:0] GEN_280;
  wire [3:0] GEN_281;
  wire  GEN_295;
  wire  GEN_296;
  wire  GEN_298;
  wire  GEN_299;
  wire  GEN_301;
  wire  GEN_302;
  wire [31:0] GEN_305;
  wire [31:0] GEN_306;
  wire  GEN_332;
  wire  GEN_333;
  wire [31:0] GEN_347;
  wire [31:0] GEN_348;
  wire [31:0] GEN_349;
  wire [31:0] GEN_350;
  wire [31:0] GEN_351;
  wire [31:0] GEN_352;
  wire  GEN_370;
  wire  GEN_371;
  wire  GEN_372;
  wire [31:0] GEN_373;
  wire [31:0] GEN_374;
  wire  GEN_378;
  wire [3:0] GEN_404;
  wire [3:0] GEN_405;
  wire  GEN_419;
  wire  GEN_420;
  wire  GEN_422;
  wire  GEN_423;
  wire  GEN_425;
  wire  GEN_426;
  wire [31:0] GEN_429;
  wire [31:0] GEN_430;
  wire  GEN_431;
  wire  GEN_432;
  wire  GEN_433;
  wire  GEN_434;
  wire  GEN_435;
  wire  GEN_436;
  reg  GEN_51;
  reg [31:0] GEN_291;
  reg [6:0] GEN_52;
  reg [31:0] GEN_292;
  reg [4:0] GEN_53;
  reg [31:0] GEN_293;
  reg [4:0] GEN_54;
  reg [31:0] GEN_294;
  reg  GEN_56;
  reg [31:0] GEN_297;
  reg  GEN_57;
  reg [31:0] GEN_300;
  reg  GEN_62;
  reg [31:0] GEN_303;
  reg [4:0] GEN_64;
  reg [31:0] GEN_304;
  reg [6:0] GEN_69;
  reg [31:0] GEN_307;
  reg [31:0] GEN_70;
  reg [31:0] GEN_308;
  reg [31:0] GEN_71;
  reg [31:0] GEN_309;
  reg  GEN_72;
  reg [31:0] GEN_310;
  reg [1:0] GEN_74;
  reg [31:0] GEN_311;
  reg  GEN_75;
  reg [31:0] GEN_312;
  reg [30:0] GEN_80;
  reg [31:0] GEN_313;
  reg  GEN_82;
  reg [31:0] GEN_314;
  reg [1:0] GEN_83;
  reg [31:0] GEN_315;
  reg [4:0] GEN_84;
  reg [31:0] GEN_316;
  reg [3:0] GEN_85;
  reg [31:0] GEN_317;
  reg  GEN_86;
  reg [31:0] GEN_318;
  reg  GEN_87;
  reg [31:0] GEN_319;
  reg  GEN_90;
  reg [31:0] GEN_320;
  reg [1:0] GEN_92;
  reg [31:0] GEN_321;
  reg [1:0] GEN_94;
  reg [31:0] GEN_322;
  reg [1:0] GEN_95;
  reg [31:0] GEN_323;
  reg [1:0] GEN_96;
  reg [31:0] GEN_324;
  reg  GEN_97;
  reg [31:0] GEN_325;
  reg  GEN_98;
  reg [31:0] GEN_326;
  reg  GEN_99;
  reg [31:0] GEN_327;
  reg  GEN_103;
  reg [31:0] GEN_328;
  reg  GEN_106;
  reg [31:0] GEN_329;
  reg  GEN_107;
  reg [31:0] GEN_330;
  reg  GEN_108;
  reg [31:0] GEN_331;
  reg  GEN_109;
  reg [31:0] GEN_334;
  reg  GEN_110;
  reg [31:0] GEN_335;
  reg  GEN_111;
  reg [31:0] GEN_336;
  reg  GEN_112;
  reg [31:0] GEN_337;
  reg  GEN_113;
  reg [31:0] GEN_338;
  reg  GEN_114;
  reg [31:0] GEN_339;
  reg [31:0] GEN_115;
  reg [31:0] GEN_340;
  reg [8:0] GEN_116;
  reg [31:0] GEN_341;
  reg [4:0] GEN_117;
  reg [31:0] GEN_342;
  reg [2:0] GEN_118;
  reg [31:0] GEN_343;
  reg [31:0] GEN_119;
  reg [31:0] GEN_344;
  reg  GEN_120;
  reg [31:0] GEN_345;
  reg  GEN_121;
  reg [31:0] GEN_346;
  reg [31:0] GEN_122;
  reg [31:0] GEN_353;
  reg [31:0] GEN_123;
  reg [31:0] GEN_354;
  reg  GEN_124;
  reg [31:0] GEN_355;
  reg  GEN_125;
  reg [31:0] GEN_356;
  reg  GEN_126;
  reg [31:0] GEN_357;
  reg  GEN_127;
  reg [31:0] GEN_358;
  reg  GEN_128;
  reg [31:0] GEN_359;
  reg  GEN_129;
  reg [31:0] GEN_360;
  reg  GEN_130;
  reg [31:0] GEN_361;
  reg  GEN_133;
  reg [31:0] GEN_362;
  reg [2:0] GEN_134;
  reg [31:0] GEN_363;
  reg  GEN_135;
  reg [31:0] GEN_364;
  reg [1:0] GEN_136;
  reg [31:0] GEN_365;
  reg  GEN_137;
  reg [31:0] GEN_366;
  reg [3:0] GEN_138;
  reg [31:0] GEN_367;
  reg [63:0] GEN_139;
  reg [63:0] GEN_368;
  reg  GEN_140;
  reg [31:0] GEN_369;
  reg  GEN_141;
  reg [31:0] GEN_375;
  reg [64:0] GEN_142;
  reg [95:0] GEN_376;
  reg [4:0] GEN_143;
  reg [31:0] GEN_377;
  reg  GEN_144;
  reg [31:0] GEN_379;
  reg  GEN_145;
  reg [31:0] GEN_380;
  assign io_rw_rdata = T_6208[31:0];
  assign io_csr_stall = reg_wfi;
  assign io_csr_xcpt = T_5991;
  assign io_eret = insn_ret;
  assign io_singleStep = T_6041;
  assign io_status_debug = reg_debug;
  assign io_status_prv = reg_mstatus_prv;
  assign io_status_sd = T_6048;
  assign io_status_zero3 = reg_mstatus_zero3;
  assign io_status_sd_rv32 = io_status_sd;
  assign io_status_zero2 = reg_mstatus_zero2;
  assign io_status_vm = reg_mstatus_vm;
  assign io_status_zero1 = reg_mstatus_zero1;
  assign io_status_mxr = reg_mstatus_mxr;
  assign io_status_pum = reg_mstatus_pum;
  assign io_status_mprv = reg_mstatus_mprv;
  assign io_status_xs = reg_mstatus_xs;
  assign io_status_fs = reg_mstatus_fs;
  assign io_status_mpp = reg_mstatus_mpp;
  assign io_status_hpp = reg_mstatus_hpp;
  assign io_status_spp = reg_mstatus_spp;
  assign io_status_mpie = reg_mstatus_mpie;
  assign io_status_hpie = reg_mstatus_hpie;
  assign io_status_spie = reg_mstatus_spie;
  assign io_status_upie = reg_mstatus_upie;
  assign io_status_mie = reg_mstatus_mie;
  assign io_status_hie = reg_mstatus_hie;
  assign io_status_sie = reg_mstatus_sie;
  assign io_status_uie = reg_mstatus_uie;
  assign io_ptbr_asid = reg_sptbr_asid;
  assign io_ptbr_ppn = reg_sptbr_ppn;
  assign io_evec = T_6038;
  assign io_fatc = insn_sfence_vm;
  assign io_time = reg_cycle[31:0];
  assign io_fcsr_rm = reg_frm;
  assign io_rocc_cmd_valid = GEN_51;
  assign io_rocc_cmd_bits_inst_funct = GEN_52;
  assign io_rocc_cmd_bits_inst_rs2 = GEN_53;
  assign io_rocc_cmd_bits_inst_rs1 = GEN_54;
  assign io_rocc_cmd_bits_inst_xd = GEN_56;
  assign io_rocc_cmd_bits_inst_xs1 = GEN_57;
  assign io_rocc_cmd_bits_inst_xs2 = GEN_62;
  assign io_rocc_cmd_bits_inst_rd = GEN_64;
  assign io_rocc_cmd_bits_inst_opcode = GEN_69;
  assign io_rocc_cmd_bits_rs1 = GEN_70;
  assign io_rocc_cmd_bits_rs2 = GEN_71;
  assign io_rocc_cmd_bits_status_debug = GEN_72;
  assign io_rocc_cmd_bits_status_prv = GEN_74;
  assign io_rocc_cmd_bits_status_sd = GEN_75;
  assign io_rocc_cmd_bits_status_zero3 = GEN_80;
  assign io_rocc_cmd_bits_status_sd_rv32 = GEN_82;
  assign io_rocc_cmd_bits_status_zero2 = GEN_83;
  assign io_rocc_cmd_bits_status_vm = GEN_84;
  assign io_rocc_cmd_bits_status_zero1 = GEN_85;
  assign io_rocc_cmd_bits_status_mxr = GEN_86;
  assign io_rocc_cmd_bits_status_pum = GEN_87;
  assign io_rocc_cmd_bits_status_mprv = GEN_90;
  assign io_rocc_cmd_bits_status_xs = GEN_92;
  assign io_rocc_cmd_bits_status_fs = GEN_94;
  assign io_rocc_cmd_bits_status_mpp = GEN_95;
  assign io_rocc_cmd_bits_status_hpp = GEN_96;
  assign io_rocc_cmd_bits_status_spp = GEN_97;
  assign io_rocc_cmd_bits_status_mpie = GEN_98;
  assign io_rocc_cmd_bits_status_hpie = GEN_99;
  assign io_rocc_cmd_bits_status_spie = GEN_103;
  assign io_rocc_cmd_bits_status_upie = GEN_106;
  assign io_rocc_cmd_bits_status_mie = GEN_107;
  assign io_rocc_cmd_bits_status_hie = GEN_108;
  assign io_rocc_cmd_bits_status_sie = GEN_109;
  assign io_rocc_cmd_bits_status_uie = GEN_110;
  assign io_rocc_resp_ready = GEN_111;
  assign io_rocc_mem_req_ready = GEN_112;
  assign io_rocc_mem_s2_nack = GEN_113;
  assign io_rocc_mem_resp_valid = GEN_114;
  assign io_rocc_mem_resp_bits_addr = GEN_115;
  assign io_rocc_mem_resp_bits_tag = GEN_116;
  assign io_rocc_mem_resp_bits_cmd = GEN_117;
  assign io_rocc_mem_resp_bits_typ = GEN_118;
  assign io_rocc_mem_resp_bits_data = GEN_119;
  assign io_rocc_mem_resp_bits_replay = GEN_120;
  assign io_rocc_mem_resp_bits_has_data = GEN_121;
  assign io_rocc_mem_resp_bits_data_word_bypass = GEN_122;
  assign io_rocc_mem_resp_bits_store_data = GEN_123;
  assign io_rocc_mem_replay_next = GEN_124;
  assign io_rocc_mem_xcpt_ma_ld = GEN_125;
  assign io_rocc_mem_xcpt_ma_st = GEN_126;
  assign io_rocc_mem_xcpt_pf_ld = GEN_127;
  assign io_rocc_mem_xcpt_pf_st = GEN_128;
  assign io_rocc_mem_ordered = GEN_129;
  assign io_rocc_autl_acquire_ready = GEN_130;
  assign io_rocc_autl_grant_valid = GEN_133;
  assign io_rocc_autl_grant_bits_addr_beat = GEN_134;
  assign io_rocc_autl_grant_bits_client_xact_id = GEN_135;
  assign io_rocc_autl_grant_bits_manager_xact_id = GEN_136;
  assign io_rocc_autl_grant_bits_is_builtin_type = GEN_137;
  assign io_rocc_autl_grant_bits_g_type = GEN_138;
  assign io_rocc_autl_grant_bits_data = GEN_139;
  assign io_rocc_fpu_req_ready = GEN_140;
  assign io_rocc_fpu_resp_valid = GEN_141;
  assign io_rocc_fpu_resp_bits_data = GEN_142;
  assign io_rocc_fpu_resp_bits_exc = GEN_143;
  assign io_rocc_exception = GEN_144;
  assign io_rocc_csr_waddr = io_rw_addr;
  assign io_rocc_csr_wdata = wdata;
  assign io_rocc_csr_wen = wen;
  assign io_rocc_host_id = GEN_145;
  assign io_interrupt = GEN_31;
  assign io_interrupt_cause = GEN_32;
  assign io_bp_0_control_tdrtype = reg_bp_0_control_tdrtype;
  assign io_bp_0_control_bpamaskmax = reg_bp_0_control_bpamaskmax;
  assign io_bp_0_control_reserved = reg_bp_0_control_reserved;
  assign io_bp_0_control_bpaction = reg_bp_0_control_bpaction;
  assign io_bp_0_control_bpmatch = reg_bp_0_control_bpmatch;
  assign io_bp_0_control_m = reg_bp_0_control_m;
  assign io_bp_0_control_h = reg_bp_0_control_h;
  assign io_bp_0_control_s = reg_bp_0_control_s;
  assign io_bp_0_control_u = reg_bp_0_control_u;
  assign io_bp_0_control_r = reg_bp_0_control_r;
  assign io_bp_0_control_w = reg_bp_0_control_w;
  assign io_bp_0_control_x = reg_bp_0_control_x;
  assign io_bp_0_address = reg_bp_0_address;
  assign io_bp_1_control_tdrtype = reg_bp_1_control_tdrtype;
  assign io_bp_1_control_bpamaskmax = reg_bp_1_control_bpamaskmax;
  assign io_bp_1_control_reserved = reg_bp_1_control_reserved;
  assign io_bp_1_control_bpaction = reg_bp_1_control_bpaction;
  assign io_bp_1_control_bpmatch = reg_bp_1_control_bpmatch;
  assign io_bp_1_control_m = reg_bp_1_control_m;
  assign io_bp_1_control_h = reg_bp_1_control_h;
  assign io_bp_1_control_s = reg_bp_1_control_s;
  assign io_bp_1_control_u = reg_bp_1_control_u;
  assign io_bp_1_control_r = reg_bp_1_control_r;
  assign io_bp_1_control_w = reg_bp_1_control_w;
  assign io_bp_1_control_x = reg_bp_1_control_x;
  assign io_bp_1_address = reg_bp_1_address;
  assign T_5012_debug = T_5062;
  assign T_5012_prv = T_5061;
  assign T_5012_sd = T_5060;
  assign T_5012_zero3 = T_5059;
  assign T_5012_sd_rv32 = T_5058;
  assign T_5012_zero2 = T_5057;
  assign T_5012_vm = T_5056;
  assign T_5012_zero1 = T_5055;
  assign T_5012_mxr = T_5054;
  assign T_5012_pum = T_5053;
  assign T_5012_mprv = T_5052;
  assign T_5012_xs = T_5051;
  assign T_5012_fs = T_5050;
  assign T_5012_mpp = T_5049;
  assign T_5012_hpp = T_5048;
  assign T_5012_spp = T_5047;
  assign T_5012_mpie = T_5046;
  assign T_5012_hpie = T_5045;
  assign T_5012_spie = T_5044;
  assign T_5012_upie = T_5043;
  assign T_5012_mie = T_5042;
  assign T_5012_hie = T_5041;
  assign T_5012_sie = T_5040;
  assign T_5012_uie = T_5039;
  assign T_5038 = 67'h0;
  assign T_5039 = T_5038[0];
  assign T_5040 = T_5038[1];
  assign T_5041 = T_5038[2];
  assign T_5042 = T_5038[3];
  assign T_5043 = T_5038[4];
  assign T_5044 = T_5038[5];
  assign T_5045 = T_5038[6];
  assign T_5046 = T_5038[7];
  assign T_5047 = T_5038[8];
  assign T_5048 = T_5038[10:9];
  assign T_5049 = T_5038[12:11];
  assign T_5050 = T_5038[14:13];
  assign T_5051 = T_5038[16:15];
  assign T_5052 = T_5038[17];
  assign T_5053 = T_5038[18];
  assign T_5054 = T_5038[19];
  assign T_5055 = T_5038[23:20];
  assign T_5056 = T_5038[28:24];
  assign T_5057 = T_5038[30:29];
  assign T_5058 = T_5038[31];
  assign T_5059 = T_5038[62:32];
  assign T_5060 = T_5038[63];
  assign T_5061 = T_5038[65:64];
  assign T_5062 = T_5038[66];
  assign reset_mstatus_debug = T_5012_debug;
  assign reset_mstatus_prv = 2'h3;
  assign reset_mstatus_sd = T_5012_sd;
  assign reset_mstatus_zero3 = T_5012_zero3;
  assign reset_mstatus_sd_rv32 = T_5012_sd_rv32;
  assign reset_mstatus_zero2 = T_5012_zero2;
  assign reset_mstatus_vm = T_5012_vm;
  assign reset_mstatus_zero1 = T_5012_zero1;
  assign reset_mstatus_mxr = T_5012_mxr;
  assign reset_mstatus_pum = T_5012_pum;
  assign reset_mstatus_mprv = T_5012_mprv;
  assign reset_mstatus_xs = T_5012_xs;
  assign reset_mstatus_fs = T_5012_fs;
  assign reset_mstatus_mpp = 2'h3;
  assign reset_mstatus_hpp = T_5012_hpp;
  assign reset_mstatus_spp = T_5012_spp;
  assign reset_mstatus_mpie = T_5012_mpie;
  assign reset_mstatus_hpie = T_5012_hpie;
  assign reset_mstatus_spie = T_5012_spie;
  assign reset_mstatus_upie = T_5012_upie;
  assign reset_mstatus_mie = T_5012_mie;
  assign reset_mstatus_hie = T_5012_hie;
  assign reset_mstatus_sie = T_5012_sie;
  assign reset_mstatus_uie = T_5012_uie;
  assign T_5150_xdebugver = T_5186;
  assign T_5150_ndreset = T_5185;
  assign T_5150_fullreset = T_5184;
  assign T_5150_hwbpcount = T_5183;
  assign T_5150_ebreakm = T_5182;
  assign T_5150_ebreakh = T_5181;
  assign T_5150_ebreaks = T_5180;
  assign T_5150_ebreaku = T_5179;
  assign T_5150_zero2 = T_5178;
  assign T_5150_stopcycle = T_5177;
  assign T_5150_stoptime = T_5176;
  assign T_5150_cause = T_5175;
  assign T_5150_debugint = T_5174;
  assign T_5150_zero1 = T_5173;
  assign T_5150_halt = T_5172;
  assign T_5150_step = T_5171;
  assign T_5150_prv = T_5170;
  assign T_5169 = 32'h0;
  assign T_5170 = T_5169[1:0];
  assign T_5171 = T_5169[2];
  assign T_5172 = T_5169[3];
  assign T_5173 = T_5169[4];
  assign T_5174 = T_5169[5];
  assign T_5175 = T_5169[8:6];
  assign T_5176 = T_5169[9];
  assign T_5177 = T_5169[10];
  assign T_5178 = T_5169[11];
  assign T_5179 = T_5169[12];
  assign T_5180 = T_5169[13];
  assign T_5181 = T_5169[14];
  assign T_5182 = T_5169[15];
  assign T_5183 = T_5169[27:16];
  assign T_5184 = T_5169[28];
  assign T_5185 = T_5169[29];
  assign T_5186 = T_5169[31:30];
  assign reset_dcsr_xdebugver = 2'h1;
  assign reset_dcsr_ndreset = T_5150_ndreset;
  assign reset_dcsr_fullreset = T_5150_fullreset;
  assign reset_dcsr_hwbpcount = T_5150_hwbpcount;
  assign reset_dcsr_ebreakm = T_5150_ebreakm;
  assign reset_dcsr_ebreakh = T_5150_ebreakh;
  assign reset_dcsr_ebreaks = T_5150_ebreaks;
  assign reset_dcsr_ebreaku = T_5150_ebreaku;
  assign reset_dcsr_zero2 = T_5150_zero2;
  assign reset_dcsr_stopcycle = T_5150_stopcycle;
  assign reset_dcsr_stoptime = T_5150_stoptime;
  assign reset_dcsr_cause = T_5150_cause;
  assign reset_dcsr_debugint = T_5150_debugint;
  assign reset_dcsr_zero1 = T_5150_zero1;
  assign reset_dcsr_halt = T_5150_halt;
  assign reset_dcsr_step = T_5150_step;
  assign reset_dcsr_prv = 2'h3;
  assign T_5252_rocc = T_5280;
  assign T_5252_meip = T_5279;
  assign T_5252_heip = T_5278;
  assign T_5252_seip = T_5277;
  assign T_5252_ueip = T_5276;
  assign T_5252_mtip = T_5275;
  assign T_5252_htip = T_5274;
  assign T_5252_stip = T_5273;
  assign T_5252_utip = T_5272;
  assign T_5252_msip = T_5271;
  assign T_5252_hsip = T_5270;
  assign T_5252_ssip = T_5269;
  assign T_5252_usip = T_5268;
  assign T_5267 = 13'h0;
  assign T_5268 = T_5267[0];
  assign T_5269 = T_5267[1];
  assign T_5270 = T_5267[2];
  assign T_5271 = T_5267[3];
  assign T_5272 = T_5267[4];
  assign T_5273 = T_5267[5];
  assign T_5274 = T_5267[6];
  assign T_5275 = T_5267[7];
  assign T_5276 = T_5267[8];
  assign T_5277 = T_5267[9];
  assign T_5278 = T_5267[10];
  assign T_5279 = T_5267[11];
  assign T_5280 = T_5267[12];
  assign T_5281_rocc = 1'h0;
  assign T_5281_meip = 1'h1;
  assign T_5281_heip = T_5252_heip;
  assign T_5281_seip = 1'h0;
  assign T_5281_ueip = T_5252_ueip;
  assign T_5281_mtip = 1'h1;
  assign T_5281_htip = T_5252_htip;
  assign T_5281_stip = 1'h0;
  assign T_5281_utip = T_5252_utip;
  assign T_5281_msip = 1'h1;
  assign T_5281_hsip = T_5252_hsip;
  assign T_5281_ssip = 1'h0;
  assign T_5281_usip = T_5252_usip;
  assign T_5302_rocc = T_5281_rocc;
  assign T_5302_meip = 1'h0;
  assign T_5302_heip = T_5281_heip;
  assign T_5302_seip = T_5281_seip;
  assign T_5302_ueip = T_5281_ueip;
  assign T_5302_mtip = 1'h0;
  assign T_5302_htip = T_5281_htip;
  assign T_5302_stip = T_5281_stip;
  assign T_5302_utip = T_5281_utip;
  assign T_5302_msip = 1'h0;
  assign T_5302_hsip = T_5281_hsip;
  assign T_5302_ssip = T_5281_ssip;
  assign T_5302_usip = T_5281_usip;
  assign T_5319 = {T_5281_hsip,T_5281_ssip};
  assign T_5320 = {T_5319,T_5281_usip};
  assign T_5321 = {T_5281_stip,T_5281_utip};
  assign T_5322 = {T_5321,T_5281_msip};
  assign T_5323 = {T_5322,T_5320};
  assign T_5324 = {T_5281_ueip,T_5281_mtip};
  assign T_5325 = {T_5324,T_5281_htip};
  assign T_5326 = {T_5281_heip,T_5281_seip};
  assign T_5327 = {T_5281_rocc,T_5281_meip};
  assign T_5328 = {T_5327,T_5326};
  assign T_5329 = {T_5328,T_5325};
  assign supported_interrupts = {T_5329,T_5323};
  assign exception = io_exception | io_csr_xcpt;
  assign T_5346 = io_retire | exception;
  assign GEN_27 = T_5346 ? 1'h1 : reg_singleStepped;
  assign T_5349 = io_singleStep == 1'h0;
  assign GEN_28 = T_5349 ? 1'h0 : GEN_27;
  assign T_5360 = reg_singleStepped == 1'h0;
  assign T_5362 = io_retire == 1'h0;
  assign T_5363 = T_5360 | T_5362;
  assign T_5364 = T_5363 | reset;
  assign T_5366 = T_5364 == 1'h0;
  assign GEN_437 = {{5'd0}, io_retire};
  assign T_5571 = T_5570 + GEN_437;
  assign T_5574 = T_5571[6];
  assign T_5576 = T_5573 + 58'h1;
  assign T_5577 = T_5576[57:0];
  assign GEN_29 = T_5574 ? T_5577 : T_5573;
  assign T_5578 = {T_5573,T_5570};
  assign T_5582 = T_5581 + 6'h1;
  assign T_5585 = T_5582[6];
  assign T_5587 = T_5584 + 58'h1;
  assign T_5588 = T_5587[57:0];
  assign GEN_30 = T_5585 ? T_5588 : T_5584;
  assign reg_cycle = {T_5584,T_5581};
  assign mip_rocc = io_rocc_interrupt;
  assign mip_meip = reg_mip_meip;
  assign mip_heip = reg_mip_heip;
  assign mip_seip = reg_mip_seip;
  assign mip_ueip = reg_mip_ueip;
  assign mip_mtip = reg_mip_mtip;
  assign mip_htip = reg_mip_htip;
  assign mip_stip = reg_mip_stip;
  assign mip_utip = reg_mip_utip;
  assign mip_msip = reg_mip_msip;
  assign mip_hsip = reg_mip_hsip;
  assign mip_ssip = reg_mip_ssip;
  assign mip_usip = reg_mip_usip;
  assign T_5602 = {mip_hsip,mip_ssip};
  assign T_5603 = {T_5602,mip_usip};
  assign T_5604 = {mip_stip,mip_utip};
  assign T_5605 = {T_5604,mip_msip};
  assign T_5606 = {T_5605,T_5603};
  assign T_5607 = {mip_ueip,mip_mtip};
  assign T_5608 = {T_5607,mip_htip};
  assign T_5609 = {mip_heip,mip_seip};
  assign T_5610 = {mip_rocc,mip_meip};
  assign T_5611 = {T_5610,T_5609};
  assign T_5612 = {T_5611,T_5608};
  assign T_5613 = {T_5612,T_5606};
  assign read_mip = T_5613 & supported_interrupts;
  assign GEN_438 = {{19'd0}, read_mip};
  assign pending_interrupts = GEN_438 & reg_mie;
  assign T_5615 = reg_debug == 1'h0;
  assign T_5617 = reg_mstatus_prv < 2'h3;
  assign T_5619 = reg_mstatus_prv == 2'h3;
  assign T_5620 = T_5619 & reg_mstatus_mie;
  assign T_5621 = T_5617 | T_5620;
  assign T_5622 = T_5615 & T_5621;
  assign T_5623 = ~ reg_mideleg;
  assign T_5624 = pending_interrupts & T_5623;
  assign m_interrupts = T_5622 ? T_5624 : 32'h0;
  assign T_5629 = reg_mstatus_prv < 2'h1;
  assign T_5631 = reg_mstatus_prv == 2'h1;
  assign T_5632 = T_5631 & reg_mstatus_sie;
  assign T_5633 = T_5629 | T_5632;
  assign T_5634 = T_5615 & T_5633;
  assign T_5635 = pending_interrupts & reg_mideleg;
  assign s_interrupts = T_5634 ? T_5635 : 32'h0;
  assign all_interrupts = m_interrupts | s_interrupts;
  assign T_5638 = all_interrupts[0];
  assign T_5639 = all_interrupts[1];
  assign T_5640 = all_interrupts[2];
  assign T_5641 = all_interrupts[3];
  assign T_5642 = all_interrupts[4];
  assign T_5643 = all_interrupts[5];
  assign T_5644 = all_interrupts[6];
  assign T_5645 = all_interrupts[7];
  assign T_5646 = all_interrupts[8];
  assign T_5647 = all_interrupts[9];
  assign T_5648 = all_interrupts[10];
  assign T_5649 = all_interrupts[11];
  assign T_5650 = all_interrupts[12];
  assign T_5651 = all_interrupts[13];
  assign T_5652 = all_interrupts[14];
  assign T_5653 = all_interrupts[15];
  assign T_5654 = all_interrupts[16];
  assign T_5655 = all_interrupts[17];
  assign T_5656 = all_interrupts[18];
  assign T_5657 = all_interrupts[19];
  assign T_5658 = all_interrupts[20];
  assign T_5659 = all_interrupts[21];
  assign T_5660 = all_interrupts[22];
  assign T_5661 = all_interrupts[23];
  assign T_5662 = all_interrupts[24];
  assign T_5663 = all_interrupts[25];
  assign T_5664 = all_interrupts[26];
  assign T_5665 = all_interrupts[27];
  assign T_5666 = all_interrupts[28];
  assign T_5667 = all_interrupts[29];
  assign T_5668 = all_interrupts[30];
  assign T_5702 = T_5668 ? 5'h1e : 5'h1f;
  assign T_5703 = T_5667 ? 5'h1d : T_5702;
  assign T_5704 = T_5666 ? 5'h1c : T_5703;
  assign T_5705 = T_5665 ? 5'h1b : T_5704;
  assign T_5706 = T_5664 ? 5'h1a : T_5705;
  assign T_5707 = T_5663 ? 5'h19 : T_5706;
  assign T_5708 = T_5662 ? 5'h18 : T_5707;
  assign T_5709 = T_5661 ? 5'h17 : T_5708;
  assign T_5710 = T_5660 ? 5'h16 : T_5709;
  assign T_5711 = T_5659 ? 5'h15 : T_5710;
  assign T_5712 = T_5658 ? 5'h14 : T_5711;
  assign T_5713 = T_5657 ? 5'h13 : T_5712;
  assign T_5714 = T_5656 ? 5'h12 : T_5713;
  assign T_5715 = T_5655 ? 5'h11 : T_5714;
  assign T_5716 = T_5654 ? 5'h10 : T_5715;
  assign T_5717 = T_5653 ? 5'hf : T_5716;
  assign T_5718 = T_5652 ? 5'he : T_5717;
  assign T_5719 = T_5651 ? 5'hd : T_5718;
  assign T_5720 = T_5650 ? 5'hc : T_5719;
  assign T_5721 = T_5649 ? 5'hb : T_5720;
  assign T_5722 = T_5648 ? 5'ha : T_5721;
  assign T_5723 = T_5647 ? 5'h9 : T_5722;
  assign T_5724 = T_5646 ? 5'h8 : T_5723;
  assign T_5725 = T_5645 ? 5'h7 : T_5724;
  assign T_5726 = T_5644 ? 5'h6 : T_5725;
  assign T_5727 = T_5643 ? 5'h5 : T_5726;
  assign T_5728 = T_5642 ? 5'h4 : T_5727;
  assign T_5729 = T_5641 ? 5'h3 : T_5728;
  assign T_5730 = T_5640 ? 5'h2 : T_5729;
  assign T_5731 = T_5639 ? 5'h1 : T_5730;
  assign T_5732 = T_5638 ? 5'h0 : T_5731;
  assign GEN_439 = {{27'd0}, T_5732};
  assign T_5733 = 32'h80000000 + GEN_439;
  assign interruptCause = T_5733[31:0];
  assign T_5735 = all_interrupts != 32'h0;
  assign T_5738 = T_5735 & T_5349;
  assign T_5739 = T_5738 | reg_singleStepped;
  assign T_5744 = reg_dcsr_debugint & T_5615;
  assign GEN_31 = T_5744 ? 1'h1 : T_5739;
  assign GEN_32 = T_5744 ? 32'h8000000d : interruptCause;
  assign system_insn = io_rw_cmd == 3'h4;
  assign T_5747 = io_rw_cmd != 3'h0;
  assign T_5749 = system_insn == 1'h0;
  assign cpu_ren = T_5747 & T_5749;
  assign T_5750 = {io_status_hie,io_status_sie};
  assign T_5751 = {T_5750,io_status_uie};
  assign T_5752 = {io_status_spie,io_status_upie};
  assign T_5753 = {T_5752,io_status_mie};
  assign T_5754 = {T_5753,T_5751};
  assign T_5755 = {io_status_spp,io_status_mpie};
  assign T_5756 = {T_5755,io_status_hpie};
  assign T_5757 = {io_status_fs,io_status_mpp};
  assign T_5758 = {T_5757,io_status_hpp};
  assign T_5759 = {T_5758,T_5756};
  assign T_5760 = {T_5759,T_5754};
  assign T_5761 = {io_status_pum,io_status_mprv};
  assign T_5762 = {T_5761,io_status_xs};
  assign T_5763 = {io_status_vm,io_status_zero1};
  assign T_5764 = {T_5763,io_status_mxr};
  assign T_5765 = {T_5764,T_5762};
  assign T_5766 = {io_status_zero3,io_status_sd_rv32};
  assign T_5767 = {T_5766,io_status_zero2};
  assign T_5768 = {io_status_debug,io_status_prv};
  assign T_5769 = {T_5768,io_status_sd};
  assign T_5770 = {T_5769,T_5767};
  assign T_5771 = {T_5770,T_5765};
  assign T_5772 = {T_5771,T_5760};
  assign read_mstatus = T_5772[31:0];
  assign T_5773 = {reg_tdrselect_tdrmode,reg_tdrselect_reserved};
  assign T_5774 = {T_5773,reg_tdrselect_tdrindex};
  assign GEN_0 = GEN_33;
  assign GEN_33 = reg_tdrselect_tdrindex ? reg_bp_1_control_r : reg_bp_0_control_r;
  assign GEN_1 = GEN_34;
  assign GEN_34 = reg_tdrselect_tdrindex ? reg_bp_1_control_w : reg_bp_0_control_w;
  assign T_5789 = {GEN_0,GEN_1};
  assign GEN_2 = GEN_35;
  assign GEN_35 = reg_tdrselect_tdrindex ? reg_bp_1_control_x : reg_bp_0_control_x;
  assign T_5790 = {T_5789,GEN_2};
  assign GEN_3 = GEN_36;
  assign GEN_36 = reg_tdrselect_tdrindex ? reg_bp_1_control_h : reg_bp_0_control_h;
  assign GEN_4 = GEN_37;
  assign GEN_37 = reg_tdrselect_tdrindex ? reg_bp_1_control_s : reg_bp_0_control_s;
  assign T_5791 = {GEN_3,GEN_4};
  assign GEN_5 = GEN_38;
  assign GEN_38 = reg_tdrselect_tdrindex ? reg_bp_1_control_u : reg_bp_0_control_u;
  assign T_5792 = {T_5791,GEN_5};
  assign T_5793 = {T_5792,T_5790};
  assign GEN_6 = GEN_39;
  assign GEN_39 = reg_tdrselect_tdrindex ? reg_bp_1_control_bpaction : reg_bp_0_control_bpaction;
  assign GEN_7 = GEN_40;
  assign GEN_40 = reg_tdrselect_tdrindex ? reg_bp_1_control_bpmatch : reg_bp_0_control_bpmatch;
  assign T_5794 = {GEN_6,GEN_7};
  assign GEN_8 = GEN_41;
  assign GEN_41 = reg_tdrselect_tdrindex ? reg_bp_1_control_m : reg_bp_0_control_m;
  assign T_5795 = {T_5794,GEN_8};
  assign GEN_9 = GEN_42;
  assign GEN_42 = reg_tdrselect_tdrindex ? reg_bp_1_control_tdrtype : reg_bp_0_control_tdrtype;
  assign GEN_10 = GEN_43;
  assign GEN_43 = reg_tdrselect_tdrindex ? reg_bp_1_control_bpamaskmax : reg_bp_0_control_bpamaskmax;
  assign T_5796 = {GEN_9,GEN_10};
  assign GEN_11 = GEN_44;
  assign GEN_44 = reg_tdrselect_tdrindex ? reg_bp_1_control_reserved : reg_bp_0_control_reserved;
  assign T_5797 = {T_5796,GEN_11};
  assign T_5798 = {T_5797,T_5795};
  assign T_5799 = {T_5798,T_5793};
  assign T_5822 = {reg_dcsr_step,reg_dcsr_prv};
  assign T_5823 = {reg_dcsr_zero1,reg_dcsr_halt};
  assign T_5824 = {T_5823,T_5822};
  assign T_5825 = {reg_dcsr_cause,reg_dcsr_debugint};
  assign T_5826 = {reg_dcsr_stopcycle,reg_dcsr_stoptime};
  assign T_5827 = {T_5826,T_5825};
  assign T_5828 = {T_5827,T_5824};
  assign T_5829 = {reg_dcsr_ebreaku,reg_dcsr_zero2};
  assign T_5830 = {reg_dcsr_ebreakh,reg_dcsr_ebreaks};
  assign T_5831 = {T_5830,T_5829};
  assign T_5832 = {reg_dcsr_hwbpcount,reg_dcsr_ebreakm};
  assign T_5833 = {reg_dcsr_xdebugver,reg_dcsr_ndreset};
  assign T_5834 = {T_5833,reg_dcsr_fullreset};
  assign T_5835 = {T_5834,T_5832};
  assign T_5836 = {T_5835,T_5831};
  assign T_5837 = {T_5836,T_5828};
  assign T_5838 = reg_cycle[63:32];
  assign T_5839 = T_5578[63:32];
  assign T_5844 = io_rw_addr == 12'h7a0;
  assign T_5846 = io_rw_addr == 12'h7a1;
  assign T_5848 = io_rw_addr == 12'h7a2;
  assign T_5850 = io_rw_addr == 12'hf13;
  assign T_5852 = io_rw_addr == 12'hf12;
  assign T_5854 = io_rw_addr == 12'hf11;
  assign T_5856 = io_rw_addr == 12'hf00;
  assign T_5858 = io_rw_addr == 12'hf02;
  assign T_5860 = io_rw_addr == 12'h310;
  assign T_5862 = io_rw_addr == 12'h701;
  assign T_5864 = io_rw_addr == 12'h700;
  assign T_5866 = io_rw_addr == 12'h702;
  assign T_5868 = io_rw_addr == 12'hf10;
  assign T_5870 = io_rw_addr == 12'h300;
  assign T_5872 = io_rw_addr == 12'h305;
  assign T_5874 = io_rw_addr == 12'h344;
  assign T_5876 = io_rw_addr == 12'h304;
  assign T_5878 = io_rw_addr == 12'h303;
  assign T_5880 = io_rw_addr == 12'h302;
  assign T_5882 = io_rw_addr == 12'h340;
  assign T_5884 = io_rw_addr == 12'h341;
  assign T_5886 = io_rw_addr == 12'h343;
  assign T_5888 = io_rw_addr == 12'h342;
  assign T_5890 = io_rw_addr == 12'hf14;
  assign T_5892 = io_rw_addr == 12'h7b0;
  assign T_5894 = io_rw_addr == 12'h7b1;
  assign T_5896 = io_rw_addr == 12'h7b2;
  assign T_5898 = io_rw_addr == 12'hf80;
  assign T_5900 = io_rw_addr == 12'hf82;
  assign T_5902 = io_rw_addr == 12'h781;
  assign T_5904 = io_rw_addr == 12'h780;
  assign T_5906 = io_rw_addr == 12'h782;
  assign T_5907 = T_5844 | T_5846;
  assign T_5908 = T_5907 | T_5848;
  assign T_5909 = T_5908 | T_5850;
  assign T_5910 = T_5909 | T_5852;
  assign T_5911 = T_5910 | T_5854;
  assign T_5912 = T_5911 | T_5856;
  assign T_5913 = T_5912 | T_5858;
  assign T_5914 = T_5913 | T_5860;
  assign T_5915 = T_5914 | T_5862;
  assign T_5916 = T_5915 | T_5864;
  assign T_5917 = T_5916 | T_5866;
  assign T_5918 = T_5917 | T_5868;
  assign T_5919 = T_5918 | T_5870;
  assign T_5920 = T_5919 | T_5872;
  assign T_5921 = T_5920 | T_5874;
  assign T_5922 = T_5921 | T_5876;
  assign T_5923 = T_5922 | T_5878;
  assign T_5924 = T_5923 | T_5880;
  assign T_5925 = T_5924 | T_5882;
  assign T_5926 = T_5925 | T_5884;
  assign T_5927 = T_5926 | T_5886;
  assign T_5928 = T_5927 | T_5888;
  assign T_5929 = T_5928 | T_5890;
  assign T_5930 = T_5929 | T_5892;
  assign T_5931 = T_5930 | T_5894;
  assign T_5932 = T_5931 | T_5896;
  assign T_5933 = T_5932 | T_5898;
  assign T_5934 = T_5933 | T_5900;
  assign T_5935 = T_5934 | T_5902;
  assign T_5936 = T_5935 | T_5904;
  assign addr_valid = T_5936 | T_5906;
  assign T_5938 = io_rw_addr[5];
  assign T_5939 = io_rw_addr[6:5];
  assign T_5940 = ~ T_5939;
  assign T_5942 = T_5940 == 2'h0;
  assign T_5943 = io_rw_addr[9:8];
  assign csr_addr_priv = {T_5942,T_5943};
  assign T_5944 = {reg_debug,reg_mstatus_prv};
  assign priv_sufficient = T_5944 >= csr_addr_priv;
  assign T_5945 = io_rw_addr[11:10];
  assign T_5946 = ~ T_5945;
  assign read_only = T_5946 == 2'h0;
  assign T_5948 = io_rw_cmd != 3'h5;
  assign T_5949 = cpu_ren & T_5948;
  assign cpu_wen = T_5949 & priv_sufficient;
  assign T_5951 = read_only == 1'h0;
  assign wen = cpu_wen & T_5951;
  assign T_5952 = io_rw_cmd == 3'h2;
  assign T_5953 = io_rw_cmd == 3'h3;
  assign T_5954 = T_5952 | T_5953;
  assign T_5956 = T_5954 ? io_rw_rdata : 32'h0;
  assign T_5957 = io_rw_cmd != 3'h3;
  assign T_5959 = T_5957 ? io_rw_wdata : 32'h0;
  assign T_5960 = T_5956 | T_5959;
  assign T_5963 = T_5953 ? io_rw_wdata : 32'h0;
  assign T_5964 = ~ T_5963;
  assign wdata = T_5960 & T_5964;
  assign do_system_insn = priv_sufficient & system_insn;
  assign T_5966 = io_rw_addr[2:0];
  assign opcode = 8'h1 << T_5966;
  assign T_5967 = opcode[0];
  assign insn_call = do_system_insn & T_5967;
  assign T_5968 = opcode[1];
  assign insn_break = do_system_insn & T_5968;
  assign T_5969 = opcode[2];
  assign insn_ret = do_system_insn & T_5969;
  assign T_5970 = opcode[4];
  assign insn_sfence_vm = do_system_insn & T_5970;
  assign T_5971 = opcode[5];
  assign insn_wfi = do_system_insn & T_5971;
  assign T_5972 = cpu_wen & read_only;
  assign T_5974 = priv_sufficient == 1'h0;
  assign T_5976 = addr_valid == 1'h0;
  assign T_5977 = T_5974 | T_5976;
  assign T_5984 = cpu_ren & T_5977;
  assign T_5985 = T_5972 | T_5984;
  assign T_5988 = system_insn & T_5974;
  assign T_5989 = T_5985 | T_5988;
  assign T_5990 = T_5989 | insn_call;
  assign T_5991 = T_5990 | insn_break;
  assign GEN_45 = insn_wfi ? 1'h1 : reg_wfi;
  assign T_5994 = pending_interrupts != 32'h0;
  assign GEN_46 = T_5994 ? 1'h0 : GEN_45;
  assign T_5997 = io_csr_xcpt == 1'h0;
  assign GEN_440 = {{2'd0}, reg_mstatus_prv};
  assign T_5999 = GEN_440 + 4'h8;
  assign T_6000 = T_5999[3:0];
  assign T_6003 = insn_break ? 2'h3 : 2'h2;
  assign T_6004 = insn_call ? T_6000 : {{2'd0}, T_6003};
  assign cause = T_5997 ? io_cause : {{28'd0}, T_6004};
  assign cause_lsbs = cause[4:0];
  assign T_6005 = cause[31];
  assign T_6007 = cause_lsbs == 5'hd;
  assign causeIsDebugInt = T_6005 & T_6007;
  assign T_6009 = cause == 32'h3;
  assign T_6010 = {reg_dcsr_ebreaks,reg_dcsr_ebreaku};
  assign T_6011 = {reg_dcsr_ebreakm,reg_dcsr_ebreakh};
  assign T_6012 = {T_6011,T_6010};
  assign T_6013 = T_6012 >> reg_mstatus_prv;
  assign T_6014 = T_6013[0];
  assign causeIsDebugBreak = T_6009 & T_6014;
  assign T_6016 = reg_singleStepped | causeIsDebugInt;
  assign T_6017 = T_6016 | causeIsDebugBreak;
  assign T_6018 = T_6017 | reg_debug;
  assign debugTVec = reg_debug ? 12'h808 : 12'h800;
  assign tvec = T_6018 ? {{20'd0}, debugTVec} : reg_mtvec;
  assign epc = T_5938 ? reg_dpc : reg_mepc;
  assign T_6038 = exception ? tvec : epc;
  assign T_6041 = reg_dcsr_step & T_5615;
  assign T_6042 = ~ io_status_fs;
  assign T_6044 = T_6042 == 2'h0;
  assign T_6045 = ~ io_status_xs;
  assign T_6047 = T_6045 == 2'h0;
  assign T_6048 = T_6044 | T_6047;
  assign T_6049 = ~ io_pc;
  assign T_6051 = T_6049 | 32'h3;
  assign T_6052 = ~ T_6051;
  assign T_6053 = read_mstatus >> reg_mstatus_prv;
  assign T_6054 = T_6053[0];
  assign T_6059 = causeIsDebugInt ? 2'h3 : 2'h1;
  assign T_6060 = reg_singleStepped ? 3'h4 : {{1'd0}, T_6059};
  assign GEN_47 = T_6018 ? 1'h1 : reg_debug;
  assign GEN_48 = T_6018 ? T_6052 : reg_dpc;
  assign GEN_49 = T_6018 ? T_6060 : reg_dcsr_cause;
  assign GEN_50 = T_6018 ? reg_mstatus_prv : reg_dcsr_prv;
  assign T_6062 = T_6018 == 1'h0;
  assign GEN_55 = {{1'd0}, reg_mstatus_spp};
  assign GEN_58 = T_6062 ? T_6052 : reg_mepc;
  assign GEN_59 = T_6062 ? cause : reg_mcause;
  assign GEN_60 = T_6062 ? io_badaddr : reg_mbadaddr;
  assign GEN_61 = T_6062 ? T_6054 : reg_mstatus_mpie;
  assign GEN_63 = T_6062 ? 1'h0 : reg_mstatus_mie;
  assign GEN_65 = exception ? GEN_47 : reg_debug;
  assign GEN_66 = exception ? GEN_48 : reg_dpc;
  assign GEN_67 = exception ? GEN_49 : reg_dcsr_cause;
  assign GEN_68 = exception ? GEN_50 : reg_dcsr_prv;
  assign GEN_73 = exception ? GEN_55 : {{1'd0}, reg_mstatus_spp};
  assign GEN_76 = exception ? GEN_58 : reg_mepc;
  assign GEN_77 = exception ? GEN_59 : reg_mcause;
  assign GEN_78 = exception ? GEN_60 : reg_mbadaddr;
  assign GEN_79 = exception ? GEN_61 : reg_mstatus_mpie;
  assign GEN_81 = exception ? GEN_63 : reg_mstatus_mie;
  assign GEN_88 = T_5938 ? 1'h0 : GEN_65;
  assign T_6088 = T_5938 == 1'h0;
  assign T_6090 = reg_mstatus_mpp[1];
  assign GEN_89 = T_6090 ? reg_mstatus_mpie : GEN_81;
  assign GEN_91 = T_6088 ? GEN_89 : GEN_81;
  assign GEN_93 = T_6088 ? 1'h0 : GEN_79;
  assign GEN_100 = insn_ret ? GEN_88 : GEN_65;
  assign GEN_101 = insn_ret ? GEN_91 : GEN_81;
  assign GEN_102 = insn_ret ? GEN_93 : GEN_79;
  assign T_6101 = {1'h0,io_csr_xcpt};
  assign GEN_441 = {{1'd0}, io_exception};
  assign T_6102 = GEN_441 + T_6101;
  assign T_6103 = T_6102[1:0];
  assign T_6104 = {1'h0,T_6103};
  assign GEN_442 = {{2'd0}, insn_ret};
  assign T_6105 = GEN_442 + T_6104;
  assign T_6106 = T_6105[2:0];
  assign T_6108 = T_6106 <= 3'h1;
  assign T_6109 = T_6108 | reset;
  assign T_6111 = T_6109 == 1'h0;
  assign T_6113 = T_5844 ? T_5774 : 32'h0;
  assign T_6115 = T_5846 ? T_5799 : 32'h0;
  assign GEN_12 = GEN_104;
  assign GEN_104 = reg_tdrselect_tdrindex ? reg_bp_1_address : reg_bp_0_address;
  assign T_6117 = T_5848 ? GEN_12 : 32'h0;
  assign T_6125 = T_5856 ? reg_cycle : 64'h0;
  assign T_6127 = T_5858 ? T_5578 : 64'h0;
  assign T_6137 = T_5868 ? 31'h40001100 : 31'h0;
  assign T_6139 = T_5870 ? read_mstatus : 32'h0;
  assign T_6141 = T_5872 ? reg_mtvec : 32'h0;
  assign T_6143 = T_5874 ? read_mip : 13'h0;
  assign T_6145 = T_5876 ? reg_mie : 32'h0;
  assign T_6147 = T_5878 ? reg_mideleg : 32'h0;
  assign T_6149 = T_5880 ? reg_medeleg : 32'h0;
  assign T_6151 = T_5882 ? reg_mscratch : 32'h0;
  assign T_6153 = T_5884 ? reg_mepc : 32'h0;
  assign T_6155 = T_5886 ? reg_mbadaddr : 32'h0;
  assign T_6157 = T_5888 ? reg_mcause : 32'h0;
  assign T_6159 = T_5890 ? io_prci_id : 1'h0;
  assign T_6161 = T_5892 ? T_5837 : 32'h0;
  assign T_6163 = T_5894 ? reg_dpc : 32'h0;
  assign T_6165 = T_5896 ? reg_dscratch : 32'h0;
  assign T_6167 = T_5898 ? T_5838 : 32'h0;
  assign T_6169 = T_5900 ? T_5839 : 32'h0;
  assign T_6177 = T_6113 | T_6115;
  assign T_6178 = T_6177 | T_6117;
  assign GEN_443 = {{32'd0}, T_6178};
  assign T_6182 = GEN_443 | T_6125;
  assign T_6183 = T_6182 | T_6127;
  assign GEN_444 = {{33'd0}, T_6137};
  assign T_6188 = T_6183 | GEN_444;
  assign GEN_445 = {{32'd0}, T_6139};
  assign T_6189 = T_6188 | GEN_445;
  assign GEN_446 = {{32'd0}, T_6141};
  assign T_6190 = T_6189 | GEN_446;
  assign GEN_447 = {{51'd0}, T_6143};
  assign T_6191 = T_6190 | GEN_447;
  assign GEN_448 = {{32'd0}, T_6145};
  assign T_6192 = T_6191 | GEN_448;
  assign GEN_449 = {{32'd0}, T_6147};
  assign T_6193 = T_6192 | GEN_449;
  assign GEN_450 = {{32'd0}, T_6149};
  assign T_6194 = T_6193 | GEN_450;
  assign GEN_451 = {{32'd0}, T_6151};
  assign T_6195 = T_6194 | GEN_451;
  assign GEN_452 = {{32'd0}, T_6153};
  assign T_6196 = T_6195 | GEN_452;
  assign GEN_453 = {{32'd0}, T_6155};
  assign T_6197 = T_6196 | GEN_453;
  assign GEN_454 = {{32'd0}, T_6157};
  assign T_6198 = T_6197 | GEN_454;
  assign GEN_455 = {{63'd0}, T_6159};
  assign T_6199 = T_6198 | GEN_455;
  assign GEN_456 = {{32'd0}, T_6161};
  assign T_6200 = T_6199 | GEN_456;
  assign GEN_457 = {{32'd0}, T_6163};
  assign T_6201 = T_6200 | GEN_457;
  assign GEN_458 = {{32'd0}, T_6165};
  assign T_6202 = T_6201 | GEN_458;
  assign GEN_459 = {{32'd0}, T_6167};
  assign T_6203 = T_6202 | GEN_459;
  assign GEN_460 = {{32'd0}, T_6169};
  assign T_6204 = T_6203 | GEN_460;
  assign T_6208 = T_6204;
  assign T_6209 = reg_fflags | io_fcsr_flags_bits;
  assign GEN_105 = io_fcsr_flags_valid ? T_6209 : reg_fflags;
  assign supportedModes_0 = 2'h3;
  assign T_6267_debug = T_6317;
  assign T_6267_prv = T_6316;
  assign T_6267_sd = T_6315;
  assign T_6267_zero3 = T_6314;
  assign T_6267_sd_rv32 = T_6313;
  assign T_6267_zero2 = T_6312;
  assign T_6267_vm = T_6311;
  assign T_6267_zero1 = T_6310;
  assign T_6267_mxr = T_6309;
  assign T_6267_pum = T_6308;
  assign T_6267_mprv = T_6307;
  assign T_6267_xs = T_6306;
  assign T_6267_fs = T_6305;
  assign T_6267_mpp = T_6304;
  assign T_6267_hpp = T_6303;
  assign T_6267_spp = T_6302;
  assign T_6267_mpie = T_6301;
  assign T_6267_hpie = T_6300;
  assign T_6267_spie = T_6299;
  assign T_6267_upie = T_6298;
  assign T_6267_mie = T_6297;
  assign T_6267_hie = T_6296;
  assign T_6267_sie = T_6295;
  assign T_6267_uie = T_6294;
  assign T_6293 = {{35'd0}, wdata};
  assign T_6294 = T_6293[0];
  assign T_6295 = T_6293[1];
  assign T_6296 = T_6293[2];
  assign T_6297 = T_6293[3];
  assign T_6298 = T_6293[4];
  assign T_6299 = T_6293[5];
  assign T_6300 = T_6293[6];
  assign T_6301 = T_6293[7];
  assign T_6302 = T_6293[8];
  assign T_6303 = T_6293[10:9];
  assign T_6304 = T_6293[12:11];
  assign T_6305 = T_6293[14:13];
  assign T_6306 = T_6293[16:15];
  assign T_6307 = T_6293[17];
  assign T_6308 = T_6293[18];
  assign T_6309 = T_6293[19];
  assign T_6310 = T_6293[23:20];
  assign T_6311 = T_6293[28:24];
  assign T_6312 = T_6293[30:29];
  assign T_6313 = T_6293[31];
  assign T_6314 = T_6293[62:32];
  assign T_6315 = T_6293[63];
  assign T_6316 = T_6293[65:64];
  assign T_6317 = T_6293[66];
  assign GEN_131 = T_5870 ? T_6267_mie : GEN_101;
  assign GEN_132 = T_5870 ? T_6267_mpie : GEN_102;
  assign T_6346_rocc = T_6372;
  assign T_6346_meip = T_6371;
  assign T_6346_heip = T_6370;
  assign T_6346_seip = T_6369;
  assign T_6346_ueip = T_6368;
  assign T_6346_mtip = T_6367;
  assign T_6346_htip = T_6366;
  assign T_6346_stip = T_6365;
  assign T_6346_utip = T_6364;
  assign T_6346_msip = T_6363;
  assign T_6346_hsip = T_6362;
  assign T_6346_ssip = T_6361;
  assign T_6346_usip = T_6360;
  assign T_6360 = wdata[0];
  assign T_6361 = wdata[1];
  assign T_6362 = wdata[2];
  assign T_6363 = wdata[3];
  assign T_6364 = wdata[4];
  assign T_6365 = wdata[5];
  assign T_6366 = wdata[6];
  assign T_6367 = wdata[7];
  assign T_6368 = wdata[8];
  assign T_6369 = wdata[9];
  assign T_6370 = wdata[10];
  assign T_6371 = wdata[11];
  assign T_6372 = wdata[12];
  assign GEN_461 = {{19'd0}, supported_interrupts};
  assign T_6373 = wdata & GEN_461;
  assign GEN_146 = T_5876 ? T_6373 : reg_mie;
  assign T_6374 = ~ wdata;
  assign T_6376 = T_6374 | 32'h3;
  assign T_6377 = ~ T_6376;
  assign GEN_147 = T_5884 ? T_6377 : GEN_76;
  assign GEN_148 = T_5882 ? wdata : reg_mscratch;
  assign T_6378 = wdata[31:2];
  assign GEN_462 = {{2'd0}, T_6378};
  assign T_6379 = GEN_462 << 2;
  assign GEN_149 = T_5872 ? T_6379 : reg_mtvec;
  assign T_6381 = wdata & 32'h8000001f;
  assign GEN_150 = T_5888 ? T_6381 : GEN_77;
  assign GEN_151 = T_5886 ? wdata : GEN_78;
  assign T_6419_xdebugver = T_6453;
  assign T_6419_ndreset = T_6452;
  assign T_6419_fullreset = T_6451;
  assign T_6419_hwbpcount = T_6450;
  assign T_6419_ebreakm = T_6449;
  assign T_6419_ebreakh = T_6448;
  assign T_6419_ebreaks = T_6447;
  assign T_6419_ebreaku = T_6372;
  assign T_6419_zero2 = T_6371;
  assign T_6419_stopcycle = T_6370;
  assign T_6419_stoptime = T_6369;
  assign T_6419_cause = T_6442;
  assign T_6419_debugint = T_6365;
  assign T_6419_zero1 = T_6364;
  assign T_6419_halt = T_6363;
  assign T_6419_step = T_6362;
  assign T_6419_prv = T_6437;
  assign T_6437 = wdata[1:0];
  assign T_6442 = wdata[8:6];
  assign T_6447 = wdata[13];
  assign T_6448 = wdata[14];
  assign T_6449 = wdata[15];
  assign T_6450 = wdata[27:16];
  assign T_6451 = wdata[28];
  assign T_6452 = wdata[29];
  assign T_6453 = wdata[31:30];
  assign GEN_169 = T_5892 ? T_6419_halt : reg_dcsr_halt;
  assign GEN_170 = T_5892 ? T_6419_step : reg_dcsr_step;
  assign GEN_171 = T_5892 ? T_6419_ebreakm : reg_dcsr_ebreakm;
  assign GEN_172 = T_5894 ? T_6377 : GEN_66;
  assign GEN_173 = T_5896 ? wdata : reg_dscratch;
  assign T_6466_tdrmode = T_6472;
  assign T_6466_reserved = T_6471;
  assign T_6466_tdrindex = T_6360;
  assign T_6471 = wdata[30:1];
  assign T_6472 = wdata[31];
  assign GEN_174 = T_5844 ? T_6466_tdrindex : reg_tdrselect_tdrindex;
  assign T_6473 = reg_tdrselect_tdrmode | reg_debug;
  assign T_6500_tdrtype = T_6524;
  assign T_6500_bpamaskmax = T_6523;
  assign T_6500_reserved = T_6522;
  assign T_6500_bpaction = T_6521;
  assign T_6500_bpmatch = T_6520;
  assign T_6500_m = T_6366;
  assign T_6500_h = T_6365;
  assign T_6500_s = T_6364;
  assign T_6500_u = T_6363;
  assign T_6500_r = T_6362;
  assign T_6500_w = T_6361;
  assign T_6500_x = T_6360;
  assign T_6520 = wdata[10:7];
  assign T_6521 = wdata[18:11];
  assign T_6522 = wdata[22:19];
  assign T_6523 = wdata[27:23];
  assign T_6524 = wdata[31:28];
  assign GEN_13 = T_6500_tdrtype;
  assign GEN_14 = T_6500_bpamaskmax;
  assign GEN_15 = T_6500_reserved;
  assign GEN_16 = T_6500_bpaction;
  assign GEN_17 = T_6500_bpmatch;
  assign GEN_183 = 1'h0 == reg_tdrselect_tdrindex ? GEN_17 : reg_bp_0_control_bpmatch;
  assign GEN_184 = reg_tdrselect_tdrindex ? GEN_17 : reg_bp_1_control_bpmatch;
  assign GEN_18 = T_6500_m;
  assign GEN_19 = T_6500_h;
  assign GEN_20 = T_6500_s;
  assign GEN_21 = T_6500_u;
  assign GEN_22 = T_6500_r;
  assign GEN_193 = 1'h0 == reg_tdrselect_tdrindex ? GEN_22 : reg_bp_0_control_r;
  assign GEN_194 = reg_tdrselect_tdrindex ? GEN_22 : reg_bp_1_control_r;
  assign GEN_23 = T_6500_w;
  assign GEN_195 = 1'h0 == reg_tdrselect_tdrindex ? GEN_23 : reg_bp_0_control_w;
  assign GEN_196 = reg_tdrselect_tdrindex ? GEN_23 : reg_bp_1_control_w;
  assign GEN_24 = T_6500_x;
  assign GEN_197 = 1'h0 == reg_tdrselect_tdrindex ? GEN_24 : reg_bp_0_control_x;
  assign GEN_198 = reg_tdrselect_tdrindex ? GEN_24 : reg_bp_1_control_x;
  assign T_6554 = T_6500_bpmatch & 4'h2;
  assign GEN_25 = T_6554;
  assign GEN_199 = 1'h0 == reg_tdrselect_tdrindex ? GEN_25 : GEN_183;
  assign GEN_200 = reg_tdrselect_tdrindex ? GEN_25 : GEN_184;
  assign GEN_226 = T_5846 ? GEN_199 : reg_bp_0_control_bpmatch;
  assign GEN_227 = T_5846 ? GEN_200 : reg_bp_1_control_bpmatch;
  assign GEN_241 = T_5846 ? GEN_193 : reg_bp_0_control_r;
  assign GEN_242 = T_5846 ? GEN_194 : reg_bp_1_control_r;
  assign GEN_244 = T_5846 ? GEN_195 : reg_bp_0_control_w;
  assign GEN_245 = T_5846 ? GEN_196 : reg_bp_1_control_w;
  assign GEN_247 = T_5846 ? GEN_197 : reg_bp_0_control_x;
  assign GEN_248 = T_5846 ? GEN_198 : reg_bp_1_control_x;
  assign GEN_26 = wdata;
  assign GEN_250 = 1'h0 == reg_tdrselect_tdrindex ? GEN_26 : reg_bp_0_address;
  assign GEN_251 = reg_tdrselect_tdrindex ? GEN_26 : reg_bp_1_address;
  assign GEN_253 = T_5848 ? GEN_250 : reg_bp_0_address;
  assign GEN_254 = T_5848 ? GEN_251 : reg_bp_1_address;
  assign GEN_280 = T_6473 ? GEN_226 : reg_bp_0_control_bpmatch;
  assign GEN_281 = T_6473 ? GEN_227 : reg_bp_1_control_bpmatch;
  assign GEN_295 = T_6473 ? GEN_241 : reg_bp_0_control_r;
  assign GEN_296 = T_6473 ? GEN_242 : reg_bp_1_control_r;
  assign GEN_298 = T_6473 ? GEN_244 : reg_bp_0_control_w;
  assign GEN_299 = T_6473 ? GEN_245 : reg_bp_1_control_w;
  assign GEN_301 = T_6473 ? GEN_247 : reg_bp_0_control_x;
  assign GEN_302 = T_6473 ? GEN_248 : reg_bp_1_control_x;
  assign GEN_305 = T_6473 ? GEN_253 : reg_bp_0_address;
  assign GEN_306 = T_6473 ? GEN_254 : reg_bp_1_address;
  assign GEN_332 = wen ? GEN_131 : GEN_101;
  assign GEN_333 = wen ? GEN_132 : GEN_102;
  assign GEN_347 = wen ? GEN_146 : reg_mie;
  assign GEN_348 = wen ? GEN_147 : GEN_76;
  assign GEN_349 = wen ? GEN_148 : reg_mscratch;
  assign GEN_350 = wen ? GEN_149 : reg_mtvec;
  assign GEN_351 = wen ? GEN_150 : GEN_77;
  assign GEN_352 = wen ? GEN_151 : GEN_78;
  assign GEN_370 = wen ? GEN_169 : reg_dcsr_halt;
  assign GEN_371 = wen ? GEN_170 : reg_dcsr_step;
  assign GEN_372 = wen ? GEN_171 : reg_dcsr_ebreakm;
  assign GEN_373 = wen ? GEN_172 : GEN_66;
  assign GEN_374 = wen ? GEN_173 : reg_dscratch;
  assign GEN_378 = wen ? GEN_174 : reg_tdrselect_tdrindex;
  assign GEN_404 = wen ? GEN_280 : reg_bp_0_control_bpmatch;
  assign GEN_405 = wen ? GEN_281 : reg_bp_1_control_bpmatch;
  assign GEN_419 = wen ? GEN_295 : reg_bp_0_control_r;
  assign GEN_420 = wen ? GEN_296 : reg_bp_1_control_r;
  assign GEN_422 = wen ? GEN_298 : reg_bp_0_control_w;
  assign GEN_423 = wen ? GEN_299 : reg_bp_1_control_w;
  assign GEN_425 = wen ? GEN_301 : reg_bp_0_control_x;
  assign GEN_426 = wen ? GEN_302 : reg_bp_1_control_x;
  assign GEN_429 = wen ? GEN_305 : reg_bp_0_address;
  assign GEN_430 = wen ? GEN_306 : reg_bp_1_address;
  assign GEN_431 = reset ? 1'h0 : GEN_419;
  assign GEN_432 = reset ? 1'h0 : GEN_422;
  assign GEN_433 = reset ? 1'h0 : GEN_425;
  assign GEN_434 = reset ? 1'h0 : GEN_420;
  assign GEN_435 = reset ? 1'h0 : GEN_423;
  assign GEN_436 = reset ? 1'h0 : GEN_426;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_152 = {1{$random}};
  reg_mstatus_debug = GEN_152[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_153 = {1{$random}};
  reg_mstatus_prv = GEN_153[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_154 = {1{$random}};
  reg_mstatus_sd = GEN_154[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_155 = {1{$random}};
  reg_mstatus_zero3 = GEN_155[30:0];
  `endif
  `ifdef RANDOMIZE
  GEN_156 = {1{$random}};
  reg_mstatus_sd_rv32 = GEN_156[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_157 = {1{$random}};
  reg_mstatus_zero2 = GEN_157[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_158 = {1{$random}};
  reg_mstatus_vm = GEN_158[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_159 = {1{$random}};
  reg_mstatus_zero1 = GEN_159[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_160 = {1{$random}};
  reg_mstatus_mxr = GEN_160[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_161 = {1{$random}};
  reg_mstatus_pum = GEN_161[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_162 = {1{$random}};
  reg_mstatus_mprv = GEN_162[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_163 = {1{$random}};
  reg_mstatus_xs = GEN_163[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_164 = {1{$random}};
  reg_mstatus_fs = GEN_164[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_165 = {1{$random}};
  reg_mstatus_mpp = GEN_165[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_166 = {1{$random}};
  reg_mstatus_hpp = GEN_166[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_167 = {1{$random}};
  reg_mstatus_spp = GEN_167[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_168 = {1{$random}};
  reg_mstatus_mpie = GEN_168[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_175 = {1{$random}};
  reg_mstatus_hpie = GEN_175[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_176 = {1{$random}};
  reg_mstatus_spie = GEN_176[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_177 = {1{$random}};
  reg_mstatus_upie = GEN_177[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_178 = {1{$random}};
  reg_mstatus_mie = GEN_178[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_179 = {1{$random}};
  reg_mstatus_hie = GEN_179[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_180 = {1{$random}};
  reg_mstatus_sie = GEN_180[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_181 = {1{$random}};
  reg_mstatus_uie = GEN_181[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_182 = {1{$random}};
  reg_dcsr_xdebugver = GEN_182[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_185 = {1{$random}};
  reg_dcsr_ndreset = GEN_185[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_186 = {1{$random}};
  reg_dcsr_fullreset = GEN_186[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_187 = {1{$random}};
  reg_dcsr_hwbpcount = GEN_187[11:0];
  `endif
  `ifdef RANDOMIZE
  GEN_188 = {1{$random}};
  reg_dcsr_ebreakm = GEN_188[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_189 = {1{$random}};
  reg_dcsr_ebreakh = GEN_189[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_190 = {1{$random}};
  reg_dcsr_ebreaks = GEN_190[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_191 = {1{$random}};
  reg_dcsr_ebreaku = GEN_191[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_192 = {1{$random}};
  reg_dcsr_zero2 = GEN_192[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_201 = {1{$random}};
  reg_dcsr_stopcycle = GEN_201[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_202 = {1{$random}};
  reg_dcsr_stoptime = GEN_202[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_203 = {1{$random}};
  reg_dcsr_cause = GEN_203[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_204 = {1{$random}};
  reg_dcsr_debugint = GEN_204[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_205 = {1{$random}};
  reg_dcsr_zero1 = GEN_205[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_206 = {1{$random}};
  reg_dcsr_halt = GEN_206[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_207 = {1{$random}};
  reg_dcsr_step = GEN_207[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_208 = {1{$random}};
  reg_dcsr_prv = GEN_208[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_209 = {1{$random}};
  reg_debug = GEN_209[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_210 = {1{$random}};
  reg_dpc = GEN_210[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_211 = {1{$random}};
  reg_dscratch = GEN_211[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_212 = {1{$random}};
  reg_singleStepped = GEN_212[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_213 = {1{$random}};
  reg_tdrselect_tdrmode = GEN_213[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_214 = {1{$random}};
  reg_tdrselect_reserved = GEN_214[29:0];
  `endif
  `ifdef RANDOMIZE
  GEN_215 = {1{$random}};
  reg_tdrselect_tdrindex = GEN_215[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_216 = {1{$random}};
  reg_bp_0_control_tdrtype = GEN_216[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_217 = {1{$random}};
  reg_bp_0_control_bpamaskmax = GEN_217[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_218 = {1{$random}};
  reg_bp_0_control_reserved = GEN_218[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_219 = {1{$random}};
  reg_bp_0_control_bpaction = GEN_219[7:0];
  `endif
  `ifdef RANDOMIZE
  GEN_220 = {1{$random}};
  reg_bp_0_control_bpmatch = GEN_220[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_221 = {1{$random}};
  reg_bp_0_control_m = GEN_221[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_222 = {1{$random}};
  reg_bp_0_control_h = GEN_222[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_223 = {1{$random}};
  reg_bp_0_control_s = GEN_223[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_224 = {1{$random}};
  reg_bp_0_control_u = GEN_224[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_225 = {1{$random}};
  reg_bp_0_control_r = GEN_225[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_228 = {1{$random}};
  reg_bp_0_control_w = GEN_228[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_229 = {1{$random}};
  reg_bp_0_control_x = GEN_229[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_230 = {1{$random}};
  reg_bp_0_address = GEN_230[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_231 = {1{$random}};
  reg_bp_1_control_tdrtype = GEN_231[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_232 = {1{$random}};
  reg_bp_1_control_bpamaskmax = GEN_232[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_233 = {1{$random}};
  reg_bp_1_control_reserved = GEN_233[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_234 = {1{$random}};
  reg_bp_1_control_bpaction = GEN_234[7:0];
  `endif
  `ifdef RANDOMIZE
  GEN_235 = {1{$random}};
  reg_bp_1_control_bpmatch = GEN_235[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_236 = {1{$random}};
  reg_bp_1_control_m = GEN_236[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_237 = {1{$random}};
  reg_bp_1_control_h = GEN_237[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_238 = {1{$random}};
  reg_bp_1_control_s = GEN_238[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_239 = {1{$random}};
  reg_bp_1_control_u = GEN_239[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_240 = {1{$random}};
  reg_bp_1_control_r = GEN_240[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_243 = {1{$random}};
  reg_bp_1_control_w = GEN_243[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_246 = {1{$random}};
  reg_bp_1_control_x = GEN_246[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_249 = {1{$random}};
  reg_bp_1_address = GEN_249[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_252 = {1{$random}};
  reg_mie = GEN_252[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_255 = {1{$random}};
  reg_mideleg = GEN_255[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_256 = {1{$random}};
  reg_medeleg = GEN_256[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_257 = {1{$random}};
  reg_mip_rocc = GEN_257[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_258 = {1{$random}};
  reg_mip_meip = GEN_258[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_259 = {1{$random}};
  reg_mip_heip = GEN_259[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_260 = {1{$random}};
  reg_mip_seip = GEN_260[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_261 = {1{$random}};
  reg_mip_ueip = GEN_261[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_262 = {1{$random}};
  reg_mip_mtip = GEN_262[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_263 = {1{$random}};
  reg_mip_htip = GEN_263[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_264 = {1{$random}};
  reg_mip_stip = GEN_264[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_265 = {1{$random}};
  reg_mip_utip = GEN_265[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_266 = {1{$random}};
  reg_mip_msip = GEN_266[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_267 = {1{$random}};
  reg_mip_hsip = GEN_267[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_268 = {1{$random}};
  reg_mip_ssip = GEN_268[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_269 = {1{$random}};
  reg_mip_usip = GEN_269[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_270 = {1{$random}};
  reg_mepc = GEN_270[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_271 = {1{$random}};
  reg_mcause = GEN_271[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_272 = {1{$random}};
  reg_mbadaddr = GEN_272[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_273 = {1{$random}};
  reg_mscratch = GEN_273[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_274 = {1{$random}};
  reg_mtvec = GEN_274[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_275 = {1{$random}};
  reg_sepc = GEN_275[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_276 = {1{$random}};
  reg_scause = GEN_276[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_277 = {1{$random}};
  reg_sbadaddr = GEN_277[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_278 = {1{$random}};
  reg_sscratch = GEN_278[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_279 = {1{$random}};
  reg_stvec = GEN_279[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_282 = {1{$random}};
  reg_sptbr_asid = GEN_282[6:0];
  `endif
  `ifdef RANDOMIZE
  GEN_283 = {1{$random}};
  reg_sptbr_ppn = GEN_283[21:0];
  `endif
  `ifdef RANDOMIZE
  GEN_284 = {1{$random}};
  reg_wfi = GEN_284[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_285 = {1{$random}};
  reg_fflags = GEN_285[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_286 = {1{$random}};
  reg_frm = GEN_286[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_287 = {1{$random}};
  T_5570 = GEN_287[5:0];
  `endif
  `ifdef RANDOMIZE
  GEN_288 = {2{$random}};
  T_5573 = GEN_288[57:0];
  `endif
  `ifdef RANDOMIZE
  GEN_289 = {1{$random}};
  T_5581 = GEN_289[5:0];
  `endif
  `ifdef RANDOMIZE
  GEN_290 = {2{$random}};
  T_5584 = GEN_290[57:0];
  `endif
  `ifdef RANDOMIZE
  GEN_291 = {1{$random}};
  GEN_51 = GEN_291[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_292 = {1{$random}};
  GEN_52 = GEN_292[6:0];
  `endif
  `ifdef RANDOMIZE
  GEN_293 = {1{$random}};
  GEN_53 = GEN_293[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_294 = {1{$random}};
  GEN_54 = GEN_294[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_297 = {1{$random}};
  GEN_56 = GEN_297[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_300 = {1{$random}};
  GEN_57 = GEN_300[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_303 = {1{$random}};
  GEN_62 = GEN_303[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_304 = {1{$random}};
  GEN_64 = GEN_304[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_307 = {1{$random}};
  GEN_69 = GEN_307[6:0];
  `endif
  `ifdef RANDOMIZE
  GEN_308 = {1{$random}};
  GEN_70 = GEN_308[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_309 = {1{$random}};
  GEN_71 = GEN_309[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_310 = {1{$random}};
  GEN_72 = GEN_310[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_311 = {1{$random}};
  GEN_74 = GEN_311[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_312 = {1{$random}};
  GEN_75 = GEN_312[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_313 = {1{$random}};
  GEN_80 = GEN_313[30:0];
  `endif
  `ifdef RANDOMIZE
  GEN_314 = {1{$random}};
  GEN_82 = GEN_314[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_315 = {1{$random}};
  GEN_83 = GEN_315[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_316 = {1{$random}};
  GEN_84 = GEN_316[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_317 = {1{$random}};
  GEN_85 = GEN_317[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_318 = {1{$random}};
  GEN_86 = GEN_318[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_319 = {1{$random}};
  GEN_87 = GEN_319[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_320 = {1{$random}};
  GEN_90 = GEN_320[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_321 = {1{$random}};
  GEN_92 = GEN_321[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_322 = {1{$random}};
  GEN_94 = GEN_322[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_323 = {1{$random}};
  GEN_95 = GEN_323[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_324 = {1{$random}};
  GEN_96 = GEN_324[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_325 = {1{$random}};
  GEN_97 = GEN_325[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_326 = {1{$random}};
  GEN_98 = GEN_326[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_327 = {1{$random}};
  GEN_99 = GEN_327[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_328 = {1{$random}};
  GEN_103 = GEN_328[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_329 = {1{$random}};
  GEN_106 = GEN_329[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_330 = {1{$random}};
  GEN_107 = GEN_330[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_331 = {1{$random}};
  GEN_108 = GEN_331[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_334 = {1{$random}};
  GEN_109 = GEN_334[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_335 = {1{$random}};
  GEN_110 = GEN_335[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_336 = {1{$random}};
  GEN_111 = GEN_336[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_337 = {1{$random}};
  GEN_112 = GEN_337[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_338 = {1{$random}};
  GEN_113 = GEN_338[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_339 = {1{$random}};
  GEN_114 = GEN_339[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_340 = {1{$random}};
  GEN_115 = GEN_340[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_341 = {1{$random}};
  GEN_116 = GEN_341[8:0];
  `endif
  `ifdef RANDOMIZE
  GEN_342 = {1{$random}};
  GEN_117 = GEN_342[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_343 = {1{$random}};
  GEN_118 = GEN_343[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_344 = {1{$random}};
  GEN_119 = GEN_344[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_345 = {1{$random}};
  GEN_120 = GEN_345[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_346 = {1{$random}};
  GEN_121 = GEN_346[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_353 = {1{$random}};
  GEN_122 = GEN_353[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_354 = {1{$random}};
  GEN_123 = GEN_354[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_355 = {1{$random}};
  GEN_124 = GEN_355[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_356 = {1{$random}};
  GEN_125 = GEN_356[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_357 = {1{$random}};
  GEN_126 = GEN_357[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_358 = {1{$random}};
  GEN_127 = GEN_358[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_359 = {1{$random}};
  GEN_128 = GEN_359[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_360 = {1{$random}};
  GEN_129 = GEN_360[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_361 = {1{$random}};
  GEN_130 = GEN_361[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_362 = {1{$random}};
  GEN_133 = GEN_362[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_363 = {1{$random}};
  GEN_134 = GEN_363[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_364 = {1{$random}};
  GEN_135 = GEN_364[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_365 = {1{$random}};
  GEN_136 = GEN_365[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_366 = {1{$random}};
  GEN_137 = GEN_366[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_367 = {1{$random}};
  GEN_138 = GEN_367[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_368 = {2{$random}};
  GEN_139 = GEN_368[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_369 = {1{$random}};
  GEN_140 = GEN_369[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_375 = {1{$random}};
  GEN_141 = GEN_375[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_376 = {3{$random}};
  GEN_142 = GEN_376[64:0];
  `endif
  `ifdef RANDOMIZE
  GEN_377 = {1{$random}};
  GEN_143 = GEN_377[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_379 = {1{$random}};
  GEN_144 = GEN_379[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_380 = {1{$random}};
  GEN_145 = GEN_380[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      reg_mstatus_debug <= reset_mstatus_debug;
    end
    if(reset) begin
      reg_mstatus_prv <= reset_mstatus_prv;
    end else begin
      reg_mstatus_prv <= 2'h3;
    end
    if(reset) begin
      reg_mstatus_sd <= reset_mstatus_sd;
    end
    if(reset) begin
      reg_mstatus_zero3 <= reset_mstatus_zero3;
    end
    if(reset) begin
      reg_mstatus_sd_rv32 <= reset_mstatus_sd_rv32;
    end
    if(reset) begin
      reg_mstatus_zero2 <= reset_mstatus_zero2;
    end
    if(reset) begin
      reg_mstatus_vm <= reset_mstatus_vm;
    end
    if(reset) begin
      reg_mstatus_zero1 <= reset_mstatus_zero1;
    end
    if(reset) begin
      reg_mstatus_mxr <= reset_mstatus_mxr;
    end
    if(reset) begin
      reg_mstatus_pum <= reset_mstatus_pum;
    end
    if(reset) begin
      reg_mstatus_mprv <= reset_mstatus_mprv;
    end else begin
      reg_mstatus_mprv <= 1'h0;
    end
    if(reset) begin
      reg_mstatus_xs <= reset_mstatus_xs;
    end
    if(reset) begin
      reg_mstatus_fs <= reset_mstatus_fs;
    end
    if(reset) begin
      reg_mstatus_mpp <= reset_mstatus_mpp;
    end else begin
      reg_mstatus_mpp <= 2'h3;
    end
    if(reset) begin
      reg_mstatus_hpp <= reset_mstatus_hpp;
    end
    if(reset) begin
      reg_mstatus_spp <= reset_mstatus_spp;
    end else begin
      reg_mstatus_spp <= GEN_73[0];
    end
    if(reset) begin
      reg_mstatus_mpie <= reset_mstatus_mpie;
    end else begin
      if(wen) begin
        if(T_5870) begin
          reg_mstatus_mpie <= T_6267_mpie;
        end else begin
          if(insn_ret) begin
            if(T_6088) begin
              reg_mstatus_mpie <= 1'h0;
            end else begin
              if(exception) begin
                if(T_6062) begin
                  reg_mstatus_mpie <= T_6054;
                end
              end
            end
          end else begin
            if(exception) begin
              if(T_6062) begin
                reg_mstatus_mpie <= T_6054;
              end
            end
          end
        end
      end else begin
        if(insn_ret) begin
          if(T_6088) begin
            reg_mstatus_mpie <= 1'h0;
          end else begin
            if(exception) begin
              if(T_6062) begin
                reg_mstatus_mpie <= T_6054;
              end
            end
          end
        end else begin
          if(exception) begin
            if(T_6062) begin
              reg_mstatus_mpie <= T_6054;
            end
          end
        end
      end
    end
    if(reset) begin
      reg_mstatus_hpie <= reset_mstatus_hpie;
    end
    if(reset) begin
      reg_mstatus_spie <= reset_mstatus_spie;
    end
    if(reset) begin
      reg_mstatus_upie <= reset_mstatus_upie;
    end
    if(reset) begin
      reg_mstatus_mie <= reset_mstatus_mie;
    end else begin
      if(wen) begin
        if(T_5870) begin
          reg_mstatus_mie <= T_6267_mie;
        end else begin
          if(insn_ret) begin
            if(T_6088) begin
              if(T_6090) begin
                reg_mstatus_mie <= reg_mstatus_mpie;
              end else begin
                if(exception) begin
                  if(T_6062) begin
                    reg_mstatus_mie <= 1'h0;
                  end
                end
              end
            end else begin
              if(exception) begin
                if(T_6062) begin
                  reg_mstatus_mie <= 1'h0;
                end
              end
            end
          end else begin
            if(exception) begin
              if(T_6062) begin
                reg_mstatus_mie <= 1'h0;
              end
            end
          end
        end
      end else begin
        if(insn_ret) begin
          if(T_6088) begin
            if(T_6090) begin
              reg_mstatus_mie <= reg_mstatus_mpie;
            end else begin
              if(exception) begin
                if(T_6062) begin
                  reg_mstatus_mie <= 1'h0;
                end
              end
            end
          end else begin
            reg_mstatus_mie <= GEN_81;
          end
        end else begin
          reg_mstatus_mie <= GEN_81;
        end
      end
    end
    if(reset) begin
      reg_mstatus_hie <= reset_mstatus_hie;
    end
    if(reset) begin
      reg_mstatus_sie <= reset_mstatus_sie;
    end
    if(reset) begin
      reg_mstatus_uie <= reset_mstatus_uie;
    end
    if(reset) begin
      reg_dcsr_xdebugver <= reset_dcsr_xdebugver;
    end
    if(reset) begin
      reg_dcsr_ndreset <= reset_dcsr_ndreset;
    end
    if(reset) begin
      reg_dcsr_fullreset <= reset_dcsr_fullreset;
    end
    if(reset) begin
      reg_dcsr_hwbpcount <= reset_dcsr_hwbpcount;
    end else begin
      reg_dcsr_hwbpcount <= 12'h2;
    end
    if(reset) begin
      reg_dcsr_ebreakm <= reset_dcsr_ebreakm;
    end else begin
      if(wen) begin
        if(T_5892) begin
          reg_dcsr_ebreakm <= T_6419_ebreakm;
        end
      end
    end
    if(reset) begin
      reg_dcsr_ebreakh <= reset_dcsr_ebreakh;
    end
    if(reset) begin
      reg_dcsr_ebreaks <= reset_dcsr_ebreaks;
    end
    if(reset) begin
      reg_dcsr_ebreaku <= reset_dcsr_ebreaku;
    end
    if(reset) begin
      reg_dcsr_zero2 <= reset_dcsr_zero2;
    end
    if(reset) begin
      reg_dcsr_stopcycle <= reset_dcsr_stopcycle;
    end
    if(reset) begin
      reg_dcsr_stoptime <= reset_dcsr_stoptime;
    end
    if(reset) begin
      reg_dcsr_cause <= reset_dcsr_cause;
    end else begin
      if(exception) begin
        if(T_6018) begin
          if(reg_singleStepped) begin
            reg_dcsr_cause <= 3'h4;
          end else begin
            reg_dcsr_cause <= {{1'd0}, T_6059};
          end
        end
      end
    end
    if(reset) begin
      reg_dcsr_debugint <= reset_dcsr_debugint;
    end else begin
      reg_dcsr_debugint <= io_prci_interrupts_debug;
    end
    if(reset) begin
      reg_dcsr_zero1 <= reset_dcsr_zero1;
    end
    if(reset) begin
      reg_dcsr_halt <= reset_dcsr_halt;
    end else begin
      if(wen) begin
        if(T_5892) begin
          reg_dcsr_halt <= T_6419_halt;
        end
      end
    end
    if(reset) begin
      reg_dcsr_step <= reset_dcsr_step;
    end else begin
      if(wen) begin
        if(T_5892) begin
          reg_dcsr_step <= T_6419_step;
        end
      end
    end
    if(reset) begin
      reg_dcsr_prv <= reset_dcsr_prv;
    end else begin
      if(exception) begin
        if(T_6018) begin
          reg_dcsr_prv <= reg_mstatus_prv;
        end
      end
    end
    if(reset) begin
      reg_debug <= 1'h0;
    end else begin
      if(insn_ret) begin
        if(T_5938) begin
          reg_debug <= 1'h0;
        end else begin
          if(exception) begin
            if(T_6018) begin
              reg_debug <= 1'h1;
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6018) begin
            reg_debug <= 1'h1;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_5894) begin
          reg_dpc <= T_6377;
        end else begin
          if(exception) begin
            if(T_6018) begin
              reg_dpc <= T_6052;
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6018) begin
            reg_dpc <= T_6052;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_5896) begin
          reg_dscratch <= wdata;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_5349) begin
        reg_singleStepped <= 1'h0;
      end else begin
        if(T_5346) begin
          reg_singleStepped <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_tdrselect_tdrmode <= 1'h1;
    end
    if(1'h0) begin
    end else begin
      reg_tdrselect_reserved <= 30'h0;
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_5844) begin
          reg_tdrselect_tdrindex <= T_6466_tdrindex;
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_tdrtype <= 4'h1;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_bpamaskmax <= 5'h4;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_reserved <= 4'h0;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_bpaction <= 8'h0;
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6473) begin
          if(T_5846) begin
            if(1'h0 == reg_tdrselect_tdrindex) begin
              reg_bp_0_control_bpmatch <= GEN_25;
            end else begin
              if(1'h0 == reg_tdrselect_tdrindex) begin
                reg_bp_0_control_bpmatch <= GEN_17;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_m <= 1'h1;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_h <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_s <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_u <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        reg_bp_0_control_r <= 1'h0;
      end else begin
        if(wen) begin
          if(T_6473) begin
            if(T_5846) begin
              if(1'h0 == reg_tdrselect_tdrindex) begin
                reg_bp_0_control_r <= GEN_22;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        reg_bp_0_control_w <= 1'h0;
      end else begin
        if(wen) begin
          if(T_6473) begin
            if(T_5846) begin
              if(1'h0 == reg_tdrselect_tdrindex) begin
                reg_bp_0_control_w <= GEN_23;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        reg_bp_0_control_x <= 1'h0;
      end else begin
        if(wen) begin
          if(T_6473) begin
            if(T_5846) begin
              if(1'h0 == reg_tdrselect_tdrindex) begin
                reg_bp_0_control_x <= GEN_24;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6473) begin
          if(T_5848) begin
            if(1'h0 == reg_tdrselect_tdrindex) begin
              reg_bp_0_address <= GEN_26;
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_tdrtype <= 4'h1;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_bpamaskmax <= 5'h4;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_reserved <= 4'h0;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_bpaction <= 8'h0;
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6473) begin
          if(T_5846) begin
            if(reg_tdrselect_tdrindex) begin
              reg_bp_1_control_bpmatch <= GEN_25;
            end else begin
              if(reg_tdrselect_tdrindex) begin
                reg_bp_1_control_bpmatch <= GEN_17;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_m <= 1'h1;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_h <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_s <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_u <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        reg_bp_1_control_r <= 1'h0;
      end else begin
        if(wen) begin
          if(T_6473) begin
            if(T_5846) begin
              if(reg_tdrselect_tdrindex) begin
                reg_bp_1_control_r <= GEN_22;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        reg_bp_1_control_w <= 1'h0;
      end else begin
        if(wen) begin
          if(T_6473) begin
            if(T_5846) begin
              if(reg_tdrselect_tdrindex) begin
                reg_bp_1_control_w <= GEN_23;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        reg_bp_1_control_x <= 1'h0;
      end else begin
        if(wen) begin
          if(T_6473) begin
            if(T_5846) begin
              if(reg_tdrselect_tdrindex) begin
                reg_bp_1_control_x <= GEN_24;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_6473) begin
          if(T_5848) begin
            if(reg_tdrselect_tdrindex) begin
              reg_bp_1_address <= GEN_26;
            end
          end
        end
      end
    end
    if(reset) begin
      reg_mie <= 32'h0;
    end else begin
      if(wen) begin
        if(T_5876) begin
          reg_mie <= T_6373;
        end
      end
    end
    if(reset) begin
      reg_mideleg <= 32'h0;
    end
    if(reset) begin
      reg_medeleg <= 32'h0;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_meip <= io_prci_interrupts_meip;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_seip <= io_prci_interrupts_seip;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_mtip <= io_prci_interrupts_mtip;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_msip <= io_prci_interrupts_msip;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_5884) begin
          reg_mepc <= T_6377;
        end else begin
          if(exception) begin
            if(T_6062) begin
              reg_mepc <= T_6052;
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6062) begin
            reg_mepc <= T_6052;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_5888) begin
          reg_mcause <= T_6381;
        end else begin
          if(exception) begin
            if(T_6062) begin
              if(T_5997) begin
                reg_mcause <= io_cause;
              end else begin
                reg_mcause <= {{28'd0}, T_6004};
              end
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6062) begin
            if(T_5997) begin
              reg_mcause <= io_cause;
            end else begin
              reg_mcause <= {{28'd0}, T_6004};
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_5886) begin
          reg_mbadaddr <= wdata;
        end else begin
          if(exception) begin
            if(T_6062) begin
              reg_mbadaddr <= io_badaddr;
            end
          end
        end
      end else begin
        if(exception) begin
          if(T_6062) begin
            reg_mbadaddr <= io_badaddr;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(wen) begin
        if(T_5882) begin
          reg_mscratch <= wdata;
        end
      end
    end
    if(reset) begin
      reg_mtvec <= 32'h1010;
    end else begin
      if(wen) begin
        if(T_5872) begin
          reg_mtvec <= T_6379;
        end
      end
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_sptbr_asid <= 7'h0;
    end
    if(1'h0) begin
    end
    if(reset) begin
      reg_wfi <= 1'h0;
    end else begin
      if(T_5994) begin
        reg_wfi <= 1'h0;
      end else begin
        if(insn_wfi) begin
          reg_wfi <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_fcsr_flags_valid) begin
        reg_fflags <= T_6209;
      end
    end
    if(1'h0) begin
    end
    if(reset) begin
      T_5570 <= 6'h0;
    end else begin
      T_5570 <= T_5571[5:0];
    end
    if(reset) begin
      T_5573 <= 58'h0;
    end else begin
      if(T_5574) begin
        T_5573 <= T_5577;
      end
    end
    if(reset) begin
      T_5581 <= 6'h0;
    end else begin
      T_5581 <= T_5582[5:0];
    end
    if(reset) begin
      T_5584 <= 58'h0;
    end else begin
      if(T_5585) begin
        T_5584 <= T_5588;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed\n    at csr.scala:185 assert(!io.singleStep || io.retire <= UInt(1))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_5366) begin
          $fwrite(32'h80000002,"Assertion failed\n    at csr.scala:186 assert(!reg_singleStepped || io.retire === UInt(0))\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_5366) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_6111) begin
          $fwrite(32'h80000002,"Assertion failed: these conditions must be mutually exclusive\n    at csr.scala:442 assert(PopCount(insn_ret :: io.exception :: io.csr_xcpt :: Nil) <= 1, ---these conditions must be mutually exclusive---)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_6111) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module BreakpointUnit(
  input   clk,
  input   reset,
  input   io_status_debug,
  input  [1:0] io_status_prv,
  input   io_status_sd,
  input  [30:0] io_status_zero3,
  input   io_status_sd_rv32,
  input  [1:0] io_status_zero2,
  input  [4:0] io_status_vm,
  input  [3:0] io_status_zero1,
  input   io_status_mxr,
  input   io_status_pum,
  input   io_status_mprv,
  input  [1:0] io_status_xs,
  input  [1:0] io_status_fs,
  input  [1:0] io_status_mpp,
  input  [1:0] io_status_hpp,
  input   io_status_spp,
  input   io_status_mpie,
  input   io_status_hpie,
  input   io_status_spie,
  input   io_status_upie,
  input   io_status_mie,
  input   io_status_hie,
  input   io_status_sie,
  input   io_status_uie,
  input  [3:0] io_bp_0_control_tdrtype,
  input  [4:0] io_bp_0_control_bpamaskmax,
  input  [3:0] io_bp_0_control_reserved,
  input  [7:0] io_bp_0_control_bpaction,
  input  [3:0] io_bp_0_control_bpmatch,
  input   io_bp_0_control_m,
  input   io_bp_0_control_h,
  input   io_bp_0_control_s,
  input   io_bp_0_control_u,
  input   io_bp_0_control_r,
  input   io_bp_0_control_w,
  input   io_bp_0_control_x,
  input  [31:0] io_bp_0_address,
  input  [3:0] io_bp_1_control_tdrtype,
  input  [4:0] io_bp_1_control_bpamaskmax,
  input  [3:0] io_bp_1_control_reserved,
  input  [7:0] io_bp_1_control_bpaction,
  input  [3:0] io_bp_1_control_bpmatch,
  input   io_bp_1_control_m,
  input   io_bp_1_control_h,
  input   io_bp_1_control_s,
  input   io_bp_1_control_u,
  input   io_bp_1_control_r,
  input   io_bp_1_control_w,
  input   io_bp_1_control_x,
  input  [31:0] io_bp_1_address,
  input  [31:0] io_pc,
  input  [31:0] io_ea,
  output  io_xcpt_if,
  output  io_xcpt_ld,
  output  io_xcpt_st
);
  wire [1:0] T_206;
  wire [1:0] T_207;
  wire [3:0] T_208;
  wire [3:0] T_209;
  wire  T_210;
  wire [31:0] T_211;
  wire  T_212;
  wire  T_214;
  wire  T_215;
  wire [1:0] T_216;
  wire  T_217;
  wire  T_218;
  wire  T_219;
  wire [2:0] T_220;
  wire  T_221;
  wire  T_222;
  wire  T_223;
  wire [3:0] T_224;
  wire [31:0] GEN_18;
  wire [31:0] T_225;
  wire [31:0] T_226;
  wire [31:0] T_240;
  wire  T_241;
  wire  T_242;
  wire [31:0] T_244;
  wire [31:0] T_258;
  wire  T_274;
  wire  T_275;
  wire  T_308;
  wire  GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire [1:0] T_310;
  wire [1:0] T_311;
  wire [3:0] T_312;
  wire [3:0] T_313;
  wire  T_314;
  wire  T_316;
  wire  T_318;
  wire  T_319;
  wire [1:0] T_320;
  wire  T_321;
  wire  T_322;
  wire  T_323;
  wire [2:0] T_324;
  wire  T_325;
  wire  T_326;
  wire  T_327;
  wire [3:0] T_328;
  wire [31:0] GEN_24;
  wire [31:0] T_329;
  wire [31:0] T_330;
  wire [31:0] T_344;
  wire  T_345;
  wire  T_346;
  wire  GEN_6;
  wire [31:0] T_362;
  wire  T_378;
  wire  T_379;
  wire  GEN_7;
  wire  T_412;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  T_420;
  wire  T_421;
  wire  T_422;
  wire  T_424;
  wire  T_425;
  wire  T_426;
  wire  T_427;
  wire  GEN_12;
  wire  T_429;
  wire  T_431;
  wire  T_432;
  wire  T_433;
  wire  T_434;
  wire  GEN_13;
  wire  T_441;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire  GEN_17;
  assign io_xcpt_if = GEN_15;
  assign io_xcpt_ld = GEN_16;
  assign io_xcpt_st = GEN_17;
  assign T_206 = {io_bp_0_control_s,io_bp_0_control_u};
  assign T_207 = {io_bp_0_control_m,io_bp_0_control_h};
  assign T_208 = {T_207,T_206};
  assign T_209 = T_208 >> io_status_prv;
  assign T_210 = T_209[0];
  assign T_211 = ~ io_pc;
  assign T_212 = io_bp_0_control_bpmatch[1];
  assign T_214 = io_bp_0_address[0];
  assign T_215 = T_212 & T_214;
  assign T_216 = {T_215,T_212};
  assign T_217 = T_216[1];
  assign T_218 = io_bp_0_address[1];
  assign T_219 = T_217 & T_218;
  assign T_220 = {T_219,T_216};
  assign T_221 = T_220[2];
  assign T_222 = io_bp_0_address[2];
  assign T_223 = T_221 & T_222;
  assign T_224 = {T_223,T_220};
  assign GEN_18 = {{28'd0}, T_224};
  assign T_225 = T_211 | GEN_18;
  assign T_226 = ~ io_bp_0_address;
  assign T_240 = T_226 | GEN_18;
  assign T_241 = T_225 == T_240;
  assign T_242 = T_241 & io_bp_0_control_x;
  assign T_244 = ~ io_ea;
  assign T_258 = T_244 | GEN_18;
  assign T_274 = T_258 == T_240;
  assign T_275 = T_274 & io_bp_0_control_r;
  assign T_308 = T_274 & io_bp_0_control_w;
  assign GEN_3 = T_210 ? T_242 : 1'h0;
  assign GEN_4 = T_210 ? T_275 : 1'h0;
  assign GEN_5 = T_210 ? T_308 : 1'h0;
  assign T_310 = {io_bp_1_control_s,io_bp_1_control_u};
  assign T_311 = {io_bp_1_control_m,io_bp_1_control_h};
  assign T_312 = {T_311,T_310};
  assign T_313 = T_312 >> io_status_prv;
  assign T_314 = T_313[0];
  assign T_316 = io_bp_1_control_bpmatch[1];
  assign T_318 = io_bp_1_address[0];
  assign T_319 = T_316 & T_318;
  assign T_320 = {T_319,T_316};
  assign T_321 = T_320[1];
  assign T_322 = io_bp_1_address[1];
  assign T_323 = T_321 & T_322;
  assign T_324 = {T_323,T_320};
  assign T_325 = T_324[2];
  assign T_326 = io_bp_1_address[2];
  assign T_327 = T_325 & T_326;
  assign T_328 = {T_327,T_324};
  assign GEN_24 = {{28'd0}, T_328};
  assign T_329 = T_211 | GEN_24;
  assign T_330 = ~ io_bp_1_address;
  assign T_344 = T_330 | GEN_24;
  assign T_345 = T_329 == T_344;
  assign T_346 = T_345 & io_bp_1_control_x;
  assign GEN_6 = T_346 ? 1'h1 : GEN_3;
  assign T_362 = T_244 | GEN_24;
  assign T_378 = T_362 == T_344;
  assign T_379 = T_378 & io_bp_1_control_r;
  assign GEN_7 = T_379 ? 1'h1 : GEN_4;
  assign T_412 = T_378 & io_bp_1_control_w;
  assign GEN_8 = T_412 ? 1'h1 : GEN_5;
  assign GEN_9 = T_314 ? GEN_6 : GEN_3;
  assign GEN_10 = T_314 ? GEN_7 : GEN_4;
  assign GEN_11 = T_314 ? GEN_8 : GEN_5;
  assign T_420 = io_bp_1_control_bpmatch == 4'h1;
  assign T_421 = T_314 & T_420;
  assign T_422 = io_pc < io_bp_0_address;
  assign T_424 = T_422 == 1'h0;
  assign T_425 = io_pc < io_bp_1_address;
  assign T_426 = T_424 & T_425;
  assign T_427 = T_426 & io_bp_1_control_x;
  assign GEN_12 = T_427 ? 1'h1 : GEN_9;
  assign T_429 = io_ea < io_bp_0_address;
  assign T_431 = T_429 == 1'h0;
  assign T_432 = io_ea < io_bp_1_address;
  assign T_433 = T_431 & T_432;
  assign T_434 = T_433 & io_bp_1_control_r;
  assign GEN_13 = T_434 ? 1'h1 : GEN_10;
  assign T_441 = T_433 & io_bp_1_control_w;
  assign GEN_14 = T_441 ? 1'h1 : GEN_11;
  assign GEN_15 = T_421 ? GEN_12 : GEN_9;
  assign GEN_16 = T_421 ? GEN_13 : GEN_10;
  assign GEN_17 = T_421 ? GEN_14 : GEN_11;
endmodule
module ALU(
  input   clk,
  input   reset,
  input   io_dw,
  input  [3:0] io_fn,
  input  [31:0] io_in2,
  input  [31:0] io_in1,
  output [31:0] io_out,
  output [31:0] io_adder_out,
  output  io_cmp_out
);
  wire  T_6;
  wire [31:0] T_7;
  wire [31:0] in2_inv;
  wire [31:0] in1_xor_in2;
  wire [32:0] T_8;
  wire [31:0] T_9;
  wire [31:0] GEN_0;
  wire [32:0] T_11;
  wire [31:0] T_12;
  wire  T_13;
  wire  T_16;
  wire  T_18;
  wire  T_19;
  wire  T_20;
  wire  T_21;
  wire  T_22;
  wire  T_23;
  wire  T_26;
  wire  T_27;
  wire  T_28;
  wire  T_29;
  wire [4:0] shamt;
  wire  T_30;
  wire  T_31;
  wire  T_32;
  wire [15:0] T_37;
  wire [31:0] T_38;
  wire [15:0] T_39;
  wire [31:0] GEN_1;
  wire [31:0] T_40;
  wire [31:0] T_42;
  wire [31:0] T_43;
  wire [23:0] T_47;
  wire [31:0] GEN_2;
  wire [31:0] T_48;
  wire [23:0] T_49;
  wire [31:0] GEN_3;
  wire [31:0] T_50;
  wire [31:0] T_52;
  wire [31:0] T_53;
  wire [27:0] T_57;
  wire [31:0] GEN_4;
  wire [31:0] T_58;
  wire [27:0] T_59;
  wire [31:0] GEN_5;
  wire [31:0] T_60;
  wire [31:0] T_62;
  wire [31:0] T_63;
  wire [29:0] T_67;
  wire [31:0] GEN_6;
  wire [31:0] T_68;
  wire [29:0] T_69;
  wire [31:0] GEN_7;
  wire [31:0] T_70;
  wire [31:0] T_72;
  wire [31:0] T_73;
  wire [30:0] T_77;
  wire [31:0] GEN_8;
  wire [31:0] T_78;
  wire [30:0] T_79;
  wire [31:0] GEN_9;
  wire [31:0] T_80;
  wire [31:0] T_82;
  wire [31:0] T_83;
  wire [31:0] shin;
  wire  T_85;
  wire  T_86;
  wire [32:0] T_87;
  wire [32:0] T_88;
  wire [32:0] T_89;
  wire [31:0] shout_r;
  wire [15:0] T_94;
  wire [31:0] T_95;
  wire [15:0] T_96;
  wire [31:0] GEN_10;
  wire [31:0] T_97;
  wire [31:0] T_99;
  wire [31:0] T_100;
  wire [23:0] T_104;
  wire [31:0] GEN_11;
  wire [31:0] T_105;
  wire [23:0] T_106;
  wire [31:0] GEN_12;
  wire [31:0] T_107;
  wire [31:0] T_109;
  wire [31:0] T_110;
  wire [27:0] T_114;
  wire [31:0] GEN_13;
  wire [31:0] T_115;
  wire [27:0] T_116;
  wire [31:0] GEN_14;
  wire [31:0] T_117;
  wire [31:0] T_119;
  wire [31:0] T_120;
  wire [29:0] T_124;
  wire [31:0] GEN_15;
  wire [31:0] T_125;
  wire [29:0] T_126;
  wire [31:0] GEN_16;
  wire [31:0] T_127;
  wire [31:0] T_129;
  wire [31:0] T_130;
  wire [30:0] T_134;
  wire [31:0] GEN_17;
  wire [31:0] T_135;
  wire [30:0] T_136;
  wire [31:0] GEN_18;
  wire [31:0] T_137;
  wire [31:0] T_139;
  wire [31:0] shout_l;
  wire [31:0] T_144;
  wire  T_145;
  wire [31:0] T_147;
  wire [31:0] shout;
  wire  T_148;
  wire  T_149;
  wire  T_150;
  wire [31:0] T_152;
  wire  T_154;
  wire  T_155;
  wire [31:0] T_156;
  wire [31:0] T_158;
  wire [31:0] logic$;
  wire  T_159;
  wire  T_160;
  wire  T_161;
  wire  T_162;
  wire  T_163;
  wire  T_164;
  wire [31:0] GEN_19;
  wire [31:0] T_165;
  wire [31:0] shift_logic;
  wire  T_166;
  wire  T_167;
  wire  T_168;
  wire [31:0] out;
  assign io_out = out;
  assign io_adder_out = T_12;
  assign io_cmp_out = T_29;
  assign T_6 = io_fn[3];
  assign T_7 = ~ io_in2;
  assign in2_inv = T_6 ? T_7 : io_in2;
  assign in1_xor_in2 = io_in1 ^ in2_inv;
  assign T_8 = io_in1 + in2_inv;
  assign T_9 = T_8[31:0];
  assign GEN_0 = {{31'd0}, T_6};
  assign T_11 = T_9 + GEN_0;
  assign T_12 = T_11[31:0];
  assign T_13 = io_fn[0];
  assign T_16 = T_6 == 1'h0;
  assign T_18 = in1_xor_in2 == 32'h0;
  assign T_19 = io_in1[31];
  assign T_20 = io_in2[31];
  assign T_21 = T_19 == T_20;
  assign T_22 = io_adder_out[31];
  assign T_23 = io_fn[1];
  assign T_26 = T_23 ? T_20 : T_19;
  assign T_27 = T_21 ? T_22 : T_26;
  assign T_28 = T_16 ? T_18 : T_27;
  assign T_29 = T_13 ^ T_28;
  assign shamt = io_in2[4:0];
  assign T_30 = io_fn == 4'h5;
  assign T_31 = io_fn == 4'hb;
  assign T_32 = T_30 | T_31;
  assign T_37 = io_in1[31:16];
  assign T_38 = {{16'd0}, T_37};
  assign T_39 = io_in1[15:0];
  assign GEN_1 = {{16'd0}, T_39};
  assign T_40 = GEN_1 << 16;
  assign T_42 = T_40 & 32'hffff0000;
  assign T_43 = T_38 | T_42;
  assign T_47 = T_43[31:8];
  assign GEN_2 = {{8'd0}, T_47};
  assign T_48 = GEN_2 & 32'hff00ff;
  assign T_49 = T_43[23:0];
  assign GEN_3 = {{8'd0}, T_49};
  assign T_50 = GEN_3 << 8;
  assign T_52 = T_50 & 32'hff00ff00;
  assign T_53 = T_48 | T_52;
  assign T_57 = T_53[31:4];
  assign GEN_4 = {{4'd0}, T_57};
  assign T_58 = GEN_4 & 32'hf0f0f0f;
  assign T_59 = T_53[27:0];
  assign GEN_5 = {{4'd0}, T_59};
  assign T_60 = GEN_5 << 4;
  assign T_62 = T_60 & 32'hf0f0f0f0;
  assign T_63 = T_58 | T_62;
  assign T_67 = T_63[31:2];
  assign GEN_6 = {{2'd0}, T_67};
  assign T_68 = GEN_6 & 32'h33333333;
  assign T_69 = T_63[29:0];
  assign GEN_7 = {{2'd0}, T_69};
  assign T_70 = GEN_7 << 2;
  assign T_72 = T_70 & 32'hcccccccc;
  assign T_73 = T_68 | T_72;
  assign T_77 = T_73[31:1];
  assign GEN_8 = {{1'd0}, T_77};
  assign T_78 = GEN_8 & 32'h55555555;
  assign T_79 = T_73[30:0];
  assign GEN_9 = {{1'd0}, T_79};
  assign T_80 = GEN_9 << 1;
  assign T_82 = T_80 & 32'haaaaaaaa;
  assign T_83 = T_78 | T_82;
  assign shin = T_32 ? io_in1 : T_83;
  assign T_85 = shin[31];
  assign T_86 = T_6 & T_85;
  assign T_87 = {T_86,shin};
  assign T_88 = $signed(T_87);
  assign T_89 = $signed(T_88) >>> shamt;
  assign shout_r = T_89[31:0];
  assign T_94 = shout_r[31:16];
  assign T_95 = {{16'd0}, T_94};
  assign T_96 = shout_r[15:0];
  assign GEN_10 = {{16'd0}, T_96};
  assign T_97 = GEN_10 << 16;
  assign T_99 = T_97 & 32'hffff0000;
  assign T_100 = T_95 | T_99;
  assign T_104 = T_100[31:8];
  assign GEN_11 = {{8'd0}, T_104};
  assign T_105 = GEN_11 & 32'hff00ff;
  assign T_106 = T_100[23:0];
  assign GEN_12 = {{8'd0}, T_106};
  assign T_107 = GEN_12 << 8;
  assign T_109 = T_107 & 32'hff00ff00;
  assign T_110 = T_105 | T_109;
  assign T_114 = T_110[31:4];
  assign GEN_13 = {{4'd0}, T_114};
  assign T_115 = GEN_13 & 32'hf0f0f0f;
  assign T_116 = T_110[27:0];
  assign GEN_14 = {{4'd0}, T_116};
  assign T_117 = GEN_14 << 4;
  assign T_119 = T_117 & 32'hf0f0f0f0;
  assign T_120 = T_115 | T_119;
  assign T_124 = T_120[31:2];
  assign GEN_15 = {{2'd0}, T_124};
  assign T_125 = GEN_15 & 32'h33333333;
  assign T_126 = T_120[29:0];
  assign GEN_16 = {{2'd0}, T_126};
  assign T_127 = GEN_16 << 2;
  assign T_129 = T_127 & 32'hcccccccc;
  assign T_130 = T_125 | T_129;
  assign T_134 = T_130[31:1];
  assign GEN_17 = {{1'd0}, T_134};
  assign T_135 = GEN_17 & 32'h55555555;
  assign T_136 = T_130[30:0];
  assign GEN_18 = {{1'd0}, T_136};
  assign T_137 = GEN_18 << 1;
  assign T_139 = T_137 & 32'haaaaaaaa;
  assign shout_l = T_135 | T_139;
  assign T_144 = T_32 ? shout_r : 32'h0;
  assign T_145 = io_fn == 4'h1;
  assign T_147 = T_145 ? shout_l : 32'h0;
  assign shout = T_144 | T_147;
  assign T_148 = io_fn == 4'h4;
  assign T_149 = io_fn == 4'h6;
  assign T_150 = T_148 | T_149;
  assign T_152 = T_150 ? in1_xor_in2 : 32'h0;
  assign T_154 = io_fn == 4'h7;
  assign T_155 = T_149 | T_154;
  assign T_156 = io_in1 & io_in2;
  assign T_158 = T_155 ? T_156 : 32'h0;
  assign logic$ = T_152 | T_158;
  assign T_159 = io_fn == 4'h2;
  assign T_160 = io_fn == 4'h3;
  assign T_161 = T_159 | T_160;
  assign T_162 = io_fn >= 4'hc;
  assign T_163 = T_161 | T_162;
  assign T_164 = T_163 & io_cmp_out;
  assign GEN_19 = {{31'd0}, T_164};
  assign T_165 = GEN_19 | logic$;
  assign shift_logic = T_165 | shout;
  assign T_166 = io_fn == 4'h0;
  assign T_167 = io_fn == 4'ha;
  assign T_168 = T_166 | T_167;
  assign out = T_168 ? io_adder_out : shift_logic;
endmodule
module MulDiv(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [3:0] io_req_bits_fn,
  input   io_req_bits_dw,
  input  [31:0] io_req_bits_in1,
  input  [31:0] io_req_bits_in2,
  input  [4:0] io_req_bits_tag,
  input   io_kill,
  input   io_resp_ready,
  output  io_resp_valid,
  output [31:0] io_resp_bits_data,
  output [4:0] io_resp_bits_tag
);
  reg [2:0] state;
  reg [31:0] GEN_14;
  reg [3:0] req_fn;
  reg [31:0] GEN_15;
  reg  req_dw;
  reg [31:0] GEN_36;
  reg [31:0] req_in1;
  reg [31:0] GEN_37;
  reg [31:0] req_in2;
  reg [31:0] GEN_38;
  reg [4:0] req_tag;
  reg [31:0] GEN_39;
  reg [5:0] count;
  reg [31:0] GEN_40;
  reg  neg_out;
  reg [31:0] GEN_41;
  reg  isMul;
  reg [31:0] GEN_42;
  reg  isHi;
  reg [31:0] GEN_43;
  reg [32:0] divisor;
  reg [63:0] GEN_44;
  reg [65:0] remainder;
  reg [95:0] GEN_45;
  wire [3:0] T_62;
  wire  T_64;
  wire [3:0] T_66;
  wire  T_68;
  wire  T_71;
  wire [3:0] T_73;
  wire  T_75;
  wire [3:0] T_77;
  wire  T_79;
  wire  T_82;
  wire  T_83;
  wire [3:0] T_85;
  wire  T_87;
  wire [3:0] T_89;
  wire  T_91;
  wire  T_94;
  wire  T_95;
  wire  T_106;
  wire  lhs_sign;
  wire [15:0] T_112;
  wire [15:0] T_114;
  wire [31:0] lhs_in;
  wire  T_122;
  wire  rhs_sign;
  wire [15:0] T_128;
  wire [15:0] T_130;
  wire [31:0] rhs_in;
  wire [32:0] T_131;
  wire [33:0] T_133;
  wire [32:0] subtractor;
  wire  less;
  wire [31:0] T_134;
  wire [32:0] T_136;
  wire [31:0] negated_remainder;
  wire  T_137;
  wire  T_138;
  wire  T_139;
  wire [65:0] GEN_0;
  wire  T_140;
  wire  T_141;
  wire [32:0] GEN_1;
  wire [65:0] GEN_2;
  wire [32:0] GEN_3;
  wire [2:0] GEN_4;
  wire  T_142;
  wire [65:0] GEN_5;
  wire [2:0] GEN_6;
  wire  T_143;
  wire [31:0] T_144;
  wire [2:0] T_145;
  wire [65:0] GEN_7;
  wire [2:0] GEN_8;
  wire  T_146;
  wire  T_147;
  wire [32:0] T_148;
  wire [64:0] T_150;
  wire [31:0] T_151;
  wire [32:0] T_152;
  wire [32:0] T_153;
  wire [32:0] T_154;
  wire [15:0] T_155;
  wire [32:0] GEN_34;
  wire [48:0] T_156;
  wire [48:0] GEN_35;
  wire [49:0] T_157;
  wire [48:0] T_158;
  wire [48:0] T_159;
  wire [15:0] T_160;
  wire [48:0] T_161;
  wire [64:0] T_162;
  wire  T_177;
  wire [32:0] T_191;
  wire [31:0] T_193;
  wire [64:0] T_194;
  wire [32:0] T_195;
  wire [31:0] T_197;
  wire [33:0] T_198;
  wire [65:0] T_199;
  wire [6:0] T_201;
  wire [5:0] T_202;
  wire  T_204;
  wire [2:0] T_206;
  wire [2:0] GEN_9;
  wire [65:0] GEN_10;
  wire [5:0] GEN_11;
  wire [2:0] GEN_12;
  wire  T_209;
  wire  T_210;
  wire  T_212;
  wire [2:0] T_214;
  wire [2:0] GEN_13;
  wire [31:0] T_218;
  wire [31:0] T_219;
  wire [31:0] T_220;
  wire  T_223;
  wire [63:0] T_224;
  wire [64:0] T_225;
  wire  T_447;
  wire  T_464;
  wire  T_467;
  wire  GEN_16;
  wire [2:0] GEN_17;
  wire [5:0] GEN_18;
  wire [65:0] GEN_19;
  wire  GEN_20;
  wire  T_469;
  wire  T_470;
  wire [2:0] GEN_21;
  wire  T_471;
  wire  T_473;
  wire  T_474;
  wire  T_475;
  wire [2:0] T_476;
  wire  T_480;
  wire  T_481;
  wire  T_482;
  wire [32:0] T_483;
  wire [2:0] GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire [5:0] GEN_25;
  wire  GEN_26;
  wire [32:0] GEN_27;
  wire [65:0] GEN_28;
  wire [3:0] GEN_29;
  wire  GEN_30;
  wire [31:0] GEN_31;
  wire [31:0] GEN_32;
  wire [4:0] GEN_33;
  wire  T_499;
  wire  T_500;
  assign io_req_ready = T_500;
  assign io_resp_valid = T_499;
  assign io_resp_bits_data = T_134;
  assign io_resp_bits_tag = req_tag;
  assign T_62 = io_req_bits_fn & 4'h4;
  assign T_64 = T_62 == 4'h0;
  assign T_66 = io_req_bits_fn & 4'h8;
  assign T_68 = T_66 == 4'h8;
  assign T_71 = T_64 | T_68;
  assign T_73 = io_req_bits_fn & 4'h5;
  assign T_75 = T_73 == 4'h1;
  assign T_77 = io_req_bits_fn & 4'h2;
  assign T_79 = T_77 == 4'h2;
  assign T_82 = T_75 | T_79;
  assign T_83 = T_82 | T_68;
  assign T_85 = io_req_bits_fn & 4'h9;
  assign T_87 = T_85 == 4'h0;
  assign T_89 = io_req_bits_fn & 4'h3;
  assign T_91 = T_89 == 4'h0;
  assign T_94 = T_87 | T_64;
  assign T_95 = T_94 | T_91;
  assign T_106 = io_req_bits_in1[31];
  assign lhs_sign = T_95 & T_106;
  assign T_112 = io_req_bits_in1[31:16];
  assign T_114 = io_req_bits_in1[15:0];
  assign lhs_in = {T_112,T_114};
  assign T_122 = io_req_bits_in2[31];
  assign rhs_sign = T_94 & T_122;
  assign T_128 = io_req_bits_in2[31:16];
  assign T_130 = io_req_bits_in2[15:0];
  assign rhs_in = {T_128,T_130};
  assign T_131 = remainder[64:32];
  assign T_133 = T_131 - divisor;
  assign subtractor = T_133[32:0];
  assign less = subtractor[32];
  assign T_134 = remainder[31:0];
  assign T_136 = 32'h0 - T_134;
  assign negated_remainder = T_136[31:0];
  assign T_137 = state == 3'h1;
  assign T_138 = remainder[31];
  assign T_139 = T_138 | isMul;
  assign GEN_0 = T_139 ? {{34'd0}, negated_remainder} : remainder;
  assign T_140 = divisor[31];
  assign T_141 = T_140 | isMul;
  assign GEN_1 = T_141 ? subtractor : divisor;
  assign GEN_2 = T_137 ? GEN_0 : remainder;
  assign GEN_3 = T_137 ? GEN_1 : divisor;
  assign GEN_4 = T_137 ? 3'h2 : state;
  assign T_142 = state == 3'h4;
  assign GEN_5 = T_142 ? {{34'd0}, negated_remainder} : GEN_2;
  assign GEN_6 = T_142 ? 3'h5 : GEN_4;
  assign T_143 = state == 3'h3;
  assign T_144 = remainder[64:33];
  assign T_145 = neg_out ? 3'h4 : 3'h5;
  assign GEN_7 = T_143 ? {{34'd0}, T_144} : GEN_5;
  assign GEN_8 = T_143 ? T_145 : GEN_6;
  assign T_146 = state == 3'h2;
  assign T_147 = T_146 & isMul;
  assign T_148 = remainder[65:33];
  assign T_150 = {T_148,T_134};
  assign T_151 = T_150[31:0];
  assign T_152 = T_150[64:32];
  assign T_153 = $signed(T_152);
  assign T_154 = $signed(divisor);
  assign T_155 = T_151[15:0];
  assign GEN_34 = {{17'd0}, T_155};
  assign T_156 = $signed(T_154) * $signed({1'b0,GEN_34});
  assign GEN_35 = {{16{T_153[32]}},T_153};
  assign T_157 = $signed(T_156) + $signed(GEN_35);
  assign T_158 = T_157[48:0];
  assign T_159 = $signed(T_158);
  assign T_160 = T_151[31:16];
  assign T_161 = $unsigned(T_159);
  assign T_162 = {T_161,T_160};
  assign T_177 = isHi == 1'h0;
  assign T_191 = T_162[64:32];
  assign T_193 = T_162[31:0];
  assign T_194 = {T_191,T_193};
  assign T_195 = T_194[64:32];
  assign T_197 = T_194[31:0];
  assign T_198 = {T_195,1'h0};
  assign T_199 = {T_198,T_197};
  assign T_201 = count + 6'h1;
  assign T_202 = T_201[5:0];
  assign T_204 = count == 6'h1;
  assign T_206 = isHi ? 3'h3 : 3'h5;
  assign GEN_9 = T_204 ? T_206 : GEN_8;
  assign GEN_10 = T_147 ? T_199 : GEN_7;
  assign GEN_11 = T_147 ? T_202 : count;
  assign GEN_12 = T_147 ? GEN_9 : GEN_8;
  assign T_209 = isMul == 1'h0;
  assign T_210 = T_146 & T_209;
  assign T_212 = count == 6'h20;
  assign T_214 = isHi ? 3'h3 : T_145;
  assign GEN_13 = T_212 ? T_214 : GEN_12;
  assign T_218 = remainder[63:32];
  assign T_219 = subtractor[31:0];
  assign T_220 = less ? T_218 : T_219;
  assign T_223 = less == 1'h0;
  assign T_224 = {T_220,T_134};
  assign T_225 = {T_224,T_223};
  assign T_447 = count == 6'h0;
  assign T_464 = T_447 & T_223;
  assign T_467 = T_464 & T_177;
  assign GEN_16 = T_467 ? 1'h0 : neg_out;
  assign GEN_17 = T_210 ? GEN_13 : GEN_12;
  assign GEN_18 = T_210 ? T_202 : GEN_11;
  assign GEN_19 = T_210 ? {{1'd0}, T_225} : GEN_10;
  assign GEN_20 = T_210 ? GEN_16 : neg_out;
  assign T_469 = io_resp_ready & io_resp_valid;
  assign T_470 = T_469 | io_kill;
  assign GEN_21 = T_470 ? 3'h0 : GEN_17;
  assign T_471 = io_req_ready & io_req_valid;
  assign T_473 = T_71 == 1'h0;
  assign T_474 = rhs_sign & T_473;
  assign T_475 = lhs_sign | T_474;
  assign T_476 = T_475 ? 3'h1 : 3'h2;
  assign T_480 = lhs_sign != rhs_sign;
  assign T_481 = T_83 ? lhs_sign : T_480;
  assign T_482 = T_473 & T_481;
  assign T_483 = {rhs_sign,rhs_in};
  assign GEN_22 = T_471 ? T_476 : GEN_21;
  assign GEN_23 = T_471 ? T_71 : isMul;
  assign GEN_24 = T_471 ? T_83 : isHi;
  assign GEN_25 = T_471 ? 6'h0 : GEN_18;
  assign GEN_26 = T_471 ? T_482 : GEN_20;
  assign GEN_27 = T_471 ? T_483 : GEN_3;
  assign GEN_28 = T_471 ? {{34'd0}, lhs_in} : GEN_19;
  assign GEN_29 = T_471 ? io_req_bits_fn : req_fn;
  assign GEN_30 = T_471 ? io_req_bits_dw : req_dw;
  assign GEN_31 = T_471 ? io_req_bits_in1 : req_in1;
  assign GEN_32 = T_471 ? io_req_bits_in2 : req_in2;
  assign GEN_33 = T_471 ? io_req_bits_tag : req_tag;
  assign T_499 = state == 3'h5;
  assign T_500 = state == 3'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_14 = {1{$random}};
  state = GEN_14[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_15 = {1{$random}};
  req_fn = GEN_15[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_36 = {1{$random}};
  req_dw = GEN_36[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_37 = {1{$random}};
  req_in1 = GEN_37[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_38 = {1{$random}};
  req_in2 = GEN_38[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_39 = {1{$random}};
  req_tag = GEN_39[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_40 = {1{$random}};
  count = GEN_40[5:0];
  `endif
  `ifdef RANDOMIZE
  GEN_41 = {1{$random}};
  neg_out = GEN_41[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_42 = {1{$random}};
  isMul = GEN_42[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_43 = {1{$random}};
  isHi = GEN_43[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_44 = {2{$random}};
  divisor = GEN_44[32:0];
  `endif
  `ifdef RANDOMIZE
  GEN_45 = {3{$random}};
  remainder = GEN_45[65:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else begin
      if(T_471) begin
        if(T_475) begin
          state <= 3'h1;
        end else begin
          state <= 3'h2;
        end
      end else begin
        if(T_470) begin
          state <= 3'h0;
        end else begin
          if(T_210) begin
            if(T_212) begin
              if(isHi) begin
                state <= 3'h3;
              end else begin
                if(neg_out) begin
                  state <= 3'h4;
                end else begin
                  state <= 3'h5;
                end
              end
            end else begin
              if(T_147) begin
                if(T_204) begin
                  if(isHi) begin
                    state <= 3'h3;
                  end else begin
                    state <= 3'h5;
                  end
                end else begin
                  if(T_143) begin
                    if(neg_out) begin
                      state <= 3'h4;
                    end else begin
                      state <= 3'h5;
                    end
                  end else begin
                    if(T_142) begin
                      state <= 3'h5;
                    end else begin
                      if(T_137) begin
                        state <= 3'h2;
                      end
                    end
                  end
                end
              end else begin
                if(T_143) begin
                  if(neg_out) begin
                    state <= 3'h4;
                  end else begin
                    state <= 3'h5;
                  end
                end else begin
                  if(T_142) begin
                    state <= 3'h5;
                  end else begin
                    if(T_137) begin
                      state <= 3'h2;
                    end
                  end
                end
              end
            end
          end else begin
            if(T_147) begin
              if(T_204) begin
                if(isHi) begin
                  state <= 3'h3;
                end else begin
                  state <= 3'h5;
                end
              end else begin
                if(T_143) begin
                  if(neg_out) begin
                    state <= 3'h4;
                  end else begin
                    state <= 3'h5;
                  end
                end else begin
                  if(T_142) begin
                    state <= 3'h5;
                  end else begin
                    if(T_137) begin
                      state <= 3'h2;
                    end
                  end
                end
              end
            end else begin
              if(T_143) begin
                state <= T_145;
              end else begin
                if(T_142) begin
                  state <= 3'h5;
                end else begin
                  if(T_137) begin
                    state <= 3'h2;
                  end
                end
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_471) begin
        req_fn <= io_req_bits_fn;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_471) begin
        req_dw <= io_req_bits_dw;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_471) begin
        req_in1 <= io_req_bits_in1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_471) begin
        req_in2 <= io_req_bits_in2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_471) begin
        req_tag <= io_req_bits_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_471) begin
        count <= 6'h0;
      end else begin
        if(T_210) begin
          count <= T_202;
        end else begin
          if(T_147) begin
            count <= T_202;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_471) begin
        neg_out <= T_482;
      end else begin
        if(T_210) begin
          if(T_467) begin
            neg_out <= 1'h0;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_471) begin
        isMul <= T_71;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_471) begin
        isHi <= T_83;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_471) begin
        divisor <= T_483;
      end else begin
        if(T_137) begin
          if(T_141) begin
            divisor <= subtractor;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_471) begin
        remainder <= {{34'd0}, lhs_in};
      end else begin
        if(T_210) begin
          remainder <= {{1'd0}, T_225};
        end else begin
          if(T_147) begin
            remainder <= T_199;
          end else begin
            if(T_143) begin
              remainder <= {{34'd0}, T_144};
            end else begin
              if(T_142) begin
                remainder <= {{34'd0}, negated_remainder};
              end else begin
                if(T_137) begin
                  if(T_139) begin
                    remainder <= {{34'd0}, negated_remainder};
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module Rocket(
  input   clk,
  input   reset,
  input   io_prci_reset,
  input   io_prci_id,
  input   io_prci_interrupts_meip,
  input   io_prci_interrupts_seip,
  input   io_prci_interrupts_debug,
  input   io_prci_interrupts_mtip,
  input   io_prci_interrupts_msip,
  output  io_imem_req_valid,
  output [31:0] io_imem_req_bits_pc,
  output  io_imem_req_bits_speculative,
  output  io_imem_resp_ready,
  input   io_imem_resp_valid,
  input  [31:0] io_imem_resp_bits_pc,
  input  [31:0] io_imem_resp_bits_data_0,
  input   io_imem_resp_bits_mask,
  input   io_imem_resp_bits_xcpt_if,
  input   io_imem_resp_bits_replay,
  input   io_imem_btb_resp_valid,
  input   io_imem_btb_resp_bits_taken,
  input   io_imem_btb_resp_bits_mask,
  input   io_imem_btb_resp_bits_bridx,
  input  [31:0] io_imem_btb_resp_bits_target,
  input   io_imem_btb_resp_bits_entry,
  input   io_imem_btb_resp_bits_bht_history,
  input  [1:0] io_imem_btb_resp_bits_bht_value,
  output  io_imem_btb_update_valid,
  output  io_imem_btb_update_bits_prediction_valid,
  output  io_imem_btb_update_bits_prediction_bits_taken,
  output  io_imem_btb_update_bits_prediction_bits_mask,
  output  io_imem_btb_update_bits_prediction_bits_bridx,
  output [31:0] io_imem_btb_update_bits_prediction_bits_target,
  output  io_imem_btb_update_bits_prediction_bits_entry,
  output  io_imem_btb_update_bits_prediction_bits_bht_history,
  output [1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
  output [31:0] io_imem_btb_update_bits_pc,
  output [31:0] io_imem_btb_update_bits_target,
  output  io_imem_btb_update_bits_taken,
  output  io_imem_btb_update_bits_isJump,
  output  io_imem_btb_update_bits_isReturn,
  output [31:0] io_imem_btb_update_bits_br_pc,
  output  io_imem_bht_update_valid,
  output  io_imem_bht_update_bits_prediction_valid,
  output  io_imem_bht_update_bits_prediction_bits_taken,
  output  io_imem_bht_update_bits_prediction_bits_mask,
  output  io_imem_bht_update_bits_prediction_bits_bridx,
  output [31:0] io_imem_bht_update_bits_prediction_bits_target,
  output  io_imem_bht_update_bits_prediction_bits_entry,
  output  io_imem_bht_update_bits_prediction_bits_bht_history,
  output [1:0] io_imem_bht_update_bits_prediction_bits_bht_value,
  output [31:0] io_imem_bht_update_bits_pc,
  output  io_imem_bht_update_bits_taken,
  output  io_imem_bht_update_bits_mispredict,
  output  io_imem_ras_update_valid,
  output  io_imem_ras_update_bits_isCall,
  output  io_imem_ras_update_bits_isReturn,
  output [31:0] io_imem_ras_update_bits_returnAddr,
  output  io_imem_ras_update_bits_prediction_valid,
  output  io_imem_ras_update_bits_prediction_bits_taken,
  output  io_imem_ras_update_bits_prediction_bits_mask,
  output  io_imem_ras_update_bits_prediction_bits_bridx,
  output [31:0] io_imem_ras_update_bits_prediction_bits_target,
  output  io_imem_ras_update_bits_prediction_bits_entry,
  output  io_imem_ras_update_bits_prediction_bits_bht_history,
  output [1:0] io_imem_ras_update_bits_prediction_bits_bht_value,
  output  io_imem_flush_icache,
  output  io_imem_flush_tlb,
  input  [31:0] io_imem_npc,
  input   io_dmem_req_ready,
  output  io_dmem_req_valid,
  output [31:0] io_dmem_req_bits_addr,
  output [8:0] io_dmem_req_bits_tag,
  output [4:0] io_dmem_req_bits_cmd,
  output [2:0] io_dmem_req_bits_typ,
  output  io_dmem_req_bits_phys,
  output [31:0] io_dmem_req_bits_data,
  output  io_dmem_s1_kill,
  output [31:0] io_dmem_s1_data,
  input   io_dmem_s2_nack,
  input   io_dmem_resp_valid,
  input  [31:0] io_dmem_resp_bits_addr,
  input  [8:0] io_dmem_resp_bits_tag,
  input  [4:0] io_dmem_resp_bits_cmd,
  input  [2:0] io_dmem_resp_bits_typ,
  input  [31:0] io_dmem_resp_bits_data,
  input   io_dmem_resp_bits_replay,
  input   io_dmem_resp_bits_has_data,
  input  [31:0] io_dmem_resp_bits_data_word_bypass,
  input  [31:0] io_dmem_resp_bits_store_data,
  input   io_dmem_replay_next,
  input   io_dmem_xcpt_ma_ld,
  input   io_dmem_xcpt_ma_st,
  input   io_dmem_xcpt_pf_ld,
  input   io_dmem_xcpt_pf_st,
  output  io_dmem_invalidate_lr,
  input   io_dmem_ordered,
  output [6:0] io_ptw_ptbr_asid,
  output [21:0] io_ptw_ptbr_ppn,
  output  io_ptw_invalidate,
  output  io_ptw_status_debug,
  output [1:0] io_ptw_status_prv,
  output  io_ptw_status_sd,
  output [30:0] io_ptw_status_zero3,
  output  io_ptw_status_sd_rv32,
  output [1:0] io_ptw_status_zero2,
  output [4:0] io_ptw_status_vm,
  output [3:0] io_ptw_status_zero1,
  output  io_ptw_status_mxr,
  output  io_ptw_status_pum,
  output  io_ptw_status_mprv,
  output [1:0] io_ptw_status_xs,
  output [1:0] io_ptw_status_fs,
  output [1:0] io_ptw_status_mpp,
  output [1:0] io_ptw_status_hpp,
  output  io_ptw_status_spp,
  output  io_ptw_status_mpie,
  output  io_ptw_status_hpie,
  output  io_ptw_status_spie,
  output  io_ptw_status_upie,
  output  io_ptw_status_mie,
  output  io_ptw_status_hie,
  output  io_ptw_status_sie,
  output  io_ptw_status_uie,
  output [31:0] io_fpu_inst,
  output [31:0] io_fpu_fromint_data,
  output [2:0] io_fpu_fcsr_rm,
  input   io_fpu_fcsr_flags_valid,
  input  [4:0] io_fpu_fcsr_flags_bits,
  input  [63:0] io_fpu_store_data,
  input  [31:0] io_fpu_toint_data,
  output  io_fpu_dmem_resp_val,
  output [2:0] io_fpu_dmem_resp_type,
  output [4:0] io_fpu_dmem_resp_tag,
  output [63:0] io_fpu_dmem_resp_data,
  output  io_fpu_valid,
  input   io_fpu_fcsr_rdy,
  input   io_fpu_nack_mem,
  input   io_fpu_illegal_rm,
  output  io_fpu_killx,
  output  io_fpu_killm,
  input  [4:0] io_fpu_dec_cmd,
  input   io_fpu_dec_ldst,
  input   io_fpu_dec_wen,
  input   io_fpu_dec_ren1,
  input   io_fpu_dec_ren2,
  input   io_fpu_dec_ren3,
  input   io_fpu_dec_swap12,
  input   io_fpu_dec_swap23,
  input   io_fpu_dec_single,
  input   io_fpu_dec_fromint,
  input   io_fpu_dec_toint,
  input   io_fpu_dec_fastpipe,
  input   io_fpu_dec_fma,
  input   io_fpu_dec_div,
  input   io_fpu_dec_sqrt,
  input   io_fpu_dec_round,
  input   io_fpu_dec_wflags,
  input   io_fpu_sboard_set,
  input   io_fpu_sboard_clr,
  input  [4:0] io_fpu_sboard_clra,
  input   io_fpu_cp_req_ready,
  output  io_fpu_cp_req_valid,
  output [4:0] io_fpu_cp_req_bits_cmd,
  output  io_fpu_cp_req_bits_ldst,
  output  io_fpu_cp_req_bits_wen,
  output  io_fpu_cp_req_bits_ren1,
  output  io_fpu_cp_req_bits_ren2,
  output  io_fpu_cp_req_bits_ren3,
  output  io_fpu_cp_req_bits_swap12,
  output  io_fpu_cp_req_bits_swap23,
  output  io_fpu_cp_req_bits_single,
  output  io_fpu_cp_req_bits_fromint,
  output  io_fpu_cp_req_bits_toint,
  output  io_fpu_cp_req_bits_fastpipe,
  output  io_fpu_cp_req_bits_fma,
  output  io_fpu_cp_req_bits_div,
  output  io_fpu_cp_req_bits_sqrt,
  output  io_fpu_cp_req_bits_round,
  output  io_fpu_cp_req_bits_wflags,
  output [2:0] io_fpu_cp_req_bits_rm,
  output [1:0] io_fpu_cp_req_bits_typ,
  output [64:0] io_fpu_cp_req_bits_in1,
  output [64:0] io_fpu_cp_req_bits_in2,
  output [64:0] io_fpu_cp_req_bits_in3,
  output  io_fpu_cp_resp_ready,
  input   io_fpu_cp_resp_valid,
  input  [64:0] io_fpu_cp_resp_bits_data,
  input  [4:0] io_fpu_cp_resp_bits_exc,
  input   io_rocc_cmd_ready,
  output  io_rocc_cmd_valid,
  output [6:0] io_rocc_cmd_bits_inst_funct,
  output [4:0] io_rocc_cmd_bits_inst_rs2,
  output [4:0] io_rocc_cmd_bits_inst_rs1,
  output  io_rocc_cmd_bits_inst_xd,
  output  io_rocc_cmd_bits_inst_xs1,
  output  io_rocc_cmd_bits_inst_xs2,
  output [4:0] io_rocc_cmd_bits_inst_rd,
  output [6:0] io_rocc_cmd_bits_inst_opcode,
  output [31:0] io_rocc_cmd_bits_rs1,
  output [31:0] io_rocc_cmd_bits_rs2,
  output  io_rocc_cmd_bits_status_debug,
  output [1:0] io_rocc_cmd_bits_status_prv,
  output  io_rocc_cmd_bits_status_sd,
  output [30:0] io_rocc_cmd_bits_status_zero3,
  output  io_rocc_cmd_bits_status_sd_rv32,
  output [1:0] io_rocc_cmd_bits_status_zero2,
  output [4:0] io_rocc_cmd_bits_status_vm,
  output [3:0] io_rocc_cmd_bits_status_zero1,
  output  io_rocc_cmd_bits_status_mxr,
  output  io_rocc_cmd_bits_status_pum,
  output  io_rocc_cmd_bits_status_mprv,
  output [1:0] io_rocc_cmd_bits_status_xs,
  output [1:0] io_rocc_cmd_bits_status_fs,
  output [1:0] io_rocc_cmd_bits_status_mpp,
  output [1:0] io_rocc_cmd_bits_status_hpp,
  output  io_rocc_cmd_bits_status_spp,
  output  io_rocc_cmd_bits_status_mpie,
  output  io_rocc_cmd_bits_status_hpie,
  output  io_rocc_cmd_bits_status_spie,
  output  io_rocc_cmd_bits_status_upie,
  output  io_rocc_cmd_bits_status_mie,
  output  io_rocc_cmd_bits_status_hie,
  output  io_rocc_cmd_bits_status_sie,
  output  io_rocc_cmd_bits_status_uie,
  output  io_rocc_resp_ready,
  input   io_rocc_resp_valid,
  input  [4:0] io_rocc_resp_bits_rd,
  input  [31:0] io_rocc_resp_bits_data,
  output  io_rocc_mem_req_ready,
  input   io_rocc_mem_req_valid,
  input  [31:0] io_rocc_mem_req_bits_addr,
  input  [8:0] io_rocc_mem_req_bits_tag,
  input  [4:0] io_rocc_mem_req_bits_cmd,
  input  [2:0] io_rocc_mem_req_bits_typ,
  input   io_rocc_mem_req_bits_phys,
  input  [31:0] io_rocc_mem_req_bits_data,
  input   io_rocc_mem_s1_kill,
  input  [31:0] io_rocc_mem_s1_data,
  output  io_rocc_mem_s2_nack,
  output  io_rocc_mem_resp_valid,
  output [31:0] io_rocc_mem_resp_bits_addr,
  output [8:0] io_rocc_mem_resp_bits_tag,
  output [4:0] io_rocc_mem_resp_bits_cmd,
  output [2:0] io_rocc_mem_resp_bits_typ,
  output [31:0] io_rocc_mem_resp_bits_data,
  output  io_rocc_mem_resp_bits_replay,
  output  io_rocc_mem_resp_bits_has_data,
  output [31:0] io_rocc_mem_resp_bits_data_word_bypass,
  output [31:0] io_rocc_mem_resp_bits_store_data,
  output  io_rocc_mem_replay_next,
  output  io_rocc_mem_xcpt_ma_ld,
  output  io_rocc_mem_xcpt_ma_st,
  output  io_rocc_mem_xcpt_pf_ld,
  output  io_rocc_mem_xcpt_pf_st,
  input   io_rocc_mem_invalidate_lr,
  output  io_rocc_mem_ordered,
  input   io_rocc_busy,
  input   io_rocc_interrupt,
  output  io_rocc_autl_acquire_ready,
  input   io_rocc_autl_acquire_valid,
  input  [25:0] io_rocc_autl_acquire_bits_addr_block,
  input   io_rocc_autl_acquire_bits_client_xact_id,
  input  [2:0] io_rocc_autl_acquire_bits_addr_beat,
  input   io_rocc_autl_acquire_bits_is_builtin_type,
  input  [2:0] io_rocc_autl_acquire_bits_a_type,
  input  [11:0] io_rocc_autl_acquire_bits_union,
  input  [63:0] io_rocc_autl_acquire_bits_data,
  input   io_rocc_autl_grant_ready,
  output  io_rocc_autl_grant_valid,
  output [2:0] io_rocc_autl_grant_bits_addr_beat,
  output  io_rocc_autl_grant_bits_client_xact_id,
  output [1:0] io_rocc_autl_grant_bits_manager_xact_id,
  output  io_rocc_autl_grant_bits_is_builtin_type,
  output [3:0] io_rocc_autl_grant_bits_g_type,
  output [63:0] io_rocc_autl_grant_bits_data,
  output  io_rocc_fpu_req_ready,
  input   io_rocc_fpu_req_valid,
  input  [4:0] io_rocc_fpu_req_bits_cmd,
  input   io_rocc_fpu_req_bits_ldst,
  input   io_rocc_fpu_req_bits_wen,
  input   io_rocc_fpu_req_bits_ren1,
  input   io_rocc_fpu_req_bits_ren2,
  input   io_rocc_fpu_req_bits_ren3,
  input   io_rocc_fpu_req_bits_swap12,
  input   io_rocc_fpu_req_bits_swap23,
  input   io_rocc_fpu_req_bits_single,
  input   io_rocc_fpu_req_bits_fromint,
  input   io_rocc_fpu_req_bits_toint,
  input   io_rocc_fpu_req_bits_fastpipe,
  input   io_rocc_fpu_req_bits_fma,
  input   io_rocc_fpu_req_bits_div,
  input   io_rocc_fpu_req_bits_sqrt,
  input   io_rocc_fpu_req_bits_round,
  input   io_rocc_fpu_req_bits_wflags,
  input  [2:0] io_rocc_fpu_req_bits_rm,
  input  [1:0] io_rocc_fpu_req_bits_typ,
  input  [64:0] io_rocc_fpu_req_bits_in1,
  input  [64:0] io_rocc_fpu_req_bits_in2,
  input  [64:0] io_rocc_fpu_req_bits_in3,
  input   io_rocc_fpu_resp_ready,
  output  io_rocc_fpu_resp_valid,
  output [64:0] io_rocc_fpu_resp_bits_data,
  output [4:0] io_rocc_fpu_resp_bits_exc,
  output  io_rocc_exception,
  output [11:0] io_rocc_csr_waddr,
  output [31:0] io_rocc_csr_wdata,
  output  io_rocc_csr_wen,
  output  io_rocc_host_id
);
  reg  ex_ctrl_legal;
  reg [31:0] GEN_271;
  reg  ex_ctrl_fp;
  reg [31:0] GEN_272;
  reg  ex_ctrl_rocc;
  reg [31:0] GEN_273;
  reg  ex_ctrl_branch;
  reg [31:0] GEN_274;
  reg  ex_ctrl_jal;
  reg [31:0] GEN_275;
  reg  ex_ctrl_jalr;
  reg [31:0] GEN_276;
  reg  ex_ctrl_rxs2;
  reg [31:0] GEN_277;
  reg  ex_ctrl_rxs1;
  reg [31:0] GEN_278;
  reg [1:0] ex_ctrl_sel_alu2;
  reg [31:0] GEN_279;
  reg [1:0] ex_ctrl_sel_alu1;
  reg [31:0] GEN_280;
  reg [2:0] ex_ctrl_sel_imm;
  reg [31:0] GEN_281;
  reg  ex_ctrl_alu_dw;
  reg [31:0] GEN_282;
  reg [3:0] ex_ctrl_alu_fn;
  reg [31:0] GEN_283;
  reg  ex_ctrl_mem;
  reg [31:0] GEN_284;
  reg [4:0] ex_ctrl_mem_cmd;
  reg [31:0] GEN_285;
  reg [2:0] ex_ctrl_mem_type;
  reg [31:0] GEN_286;
  reg  ex_ctrl_rfs1;
  reg [31:0] GEN_287;
  reg  ex_ctrl_rfs2;
  reg [31:0] GEN_288;
  reg  ex_ctrl_rfs3;
  reg [31:0] GEN_289;
  reg  ex_ctrl_wfd;
  reg [31:0] GEN_290;
  reg  ex_ctrl_div;
  reg [31:0] GEN_291;
  reg  ex_ctrl_wxd;
  reg [31:0] GEN_292;
  reg [2:0] ex_ctrl_csr;
  reg [31:0] GEN_293;
  reg  ex_ctrl_fence_i;
  reg [31:0] GEN_294;
  reg  ex_ctrl_fence;
  reg [31:0] GEN_295;
  reg  ex_ctrl_amo;
  reg [31:0] GEN_296;
  reg  mem_ctrl_legal;
  reg [31:0] GEN_297;
  reg  mem_ctrl_fp;
  reg [31:0] GEN_298;
  reg  mem_ctrl_rocc;
  reg [31:0] GEN_299;
  reg  mem_ctrl_branch;
  reg [31:0] GEN_300;
  reg  mem_ctrl_jal;
  reg [31:0] GEN_301;
  reg  mem_ctrl_jalr;
  reg [31:0] GEN_302;
  reg  mem_ctrl_rxs2;
  reg [31:0] GEN_303;
  reg  mem_ctrl_rxs1;
  reg [31:0] GEN_304;
  reg [1:0] mem_ctrl_sel_alu2;
  reg [31:0] GEN_305;
  reg [1:0] mem_ctrl_sel_alu1;
  reg [31:0] GEN_306;
  reg [2:0] mem_ctrl_sel_imm;
  reg [31:0] GEN_307;
  reg  mem_ctrl_alu_dw;
  reg [31:0] GEN_308;
  reg [3:0] mem_ctrl_alu_fn;
  reg [31:0] GEN_309;
  reg  mem_ctrl_mem;
  reg [31:0] GEN_310;
  reg [4:0] mem_ctrl_mem_cmd;
  reg [31:0] GEN_311;
  reg [2:0] mem_ctrl_mem_type;
  reg [31:0] GEN_312;
  reg  mem_ctrl_rfs1;
  reg [31:0] GEN_313;
  reg  mem_ctrl_rfs2;
  reg [31:0] GEN_314;
  reg  mem_ctrl_rfs3;
  reg [31:0] GEN_315;
  reg  mem_ctrl_wfd;
  reg [31:0] GEN_316;
  reg  mem_ctrl_div;
  reg [31:0] GEN_317;
  reg  mem_ctrl_wxd;
  reg [31:0] GEN_318;
  reg [2:0] mem_ctrl_csr;
  reg [31:0] GEN_319;
  reg  mem_ctrl_fence_i;
  reg [31:0] GEN_320;
  reg  mem_ctrl_fence;
  reg [31:0] GEN_321;
  reg  mem_ctrl_amo;
  reg [31:0] GEN_322;
  reg  wb_ctrl_legal;
  reg [31:0] GEN_323;
  reg  wb_ctrl_fp;
  reg [31:0] GEN_324;
  reg  wb_ctrl_rocc;
  reg [31:0] GEN_325;
  reg  wb_ctrl_branch;
  reg [31:0] GEN_326;
  reg  wb_ctrl_jal;
  reg [31:0] GEN_327;
  reg  wb_ctrl_jalr;
  reg [31:0] GEN_328;
  reg  wb_ctrl_rxs2;
  reg [31:0] GEN_329;
  reg  wb_ctrl_rxs1;
  reg [31:0] GEN_330;
  reg [1:0] wb_ctrl_sel_alu2;
  reg [31:0] GEN_331;
  reg [1:0] wb_ctrl_sel_alu1;
  reg [31:0] GEN_332;
  reg [2:0] wb_ctrl_sel_imm;
  reg [31:0] GEN_333;
  reg  wb_ctrl_alu_dw;
  reg [31:0] GEN_334;
  reg [3:0] wb_ctrl_alu_fn;
  reg [31:0] GEN_335;
  reg  wb_ctrl_mem;
  reg [31:0] GEN_336;
  reg [4:0] wb_ctrl_mem_cmd;
  reg [31:0] GEN_337;
  reg [2:0] wb_ctrl_mem_type;
  reg [31:0] GEN_338;
  reg  wb_ctrl_rfs1;
  reg [31:0] GEN_339;
  reg  wb_ctrl_rfs2;
  reg [31:0] GEN_340;
  reg  wb_ctrl_rfs3;
  reg [31:0] GEN_341;
  reg  wb_ctrl_wfd;
  reg [31:0] GEN_342;
  reg  wb_ctrl_div;
  reg [31:0] GEN_343;
  reg  wb_ctrl_wxd;
  reg [31:0] GEN_344;
  reg [2:0] wb_ctrl_csr;
  reg [31:0] GEN_345;
  reg  wb_ctrl_fence_i;
  reg [31:0] GEN_346;
  reg  wb_ctrl_fence;
  reg [31:0] GEN_347;
  reg  wb_ctrl_amo;
  reg [31:0] GEN_348;
  reg  ex_reg_xcpt_interrupt;
  reg [31:0] GEN_349;
  reg  ex_reg_valid;
  reg [31:0] GEN_350;
  reg  ex_reg_btb_hit;
  reg [31:0] GEN_351;
  reg  ex_reg_btb_resp_taken;
  reg [31:0] GEN_352;
  reg  ex_reg_btb_resp_mask;
  reg [31:0] GEN_353;
  reg  ex_reg_btb_resp_bridx;
  reg [31:0] GEN_354;
  reg [31:0] ex_reg_btb_resp_target;
  reg [31:0] GEN_355;
  reg  ex_reg_btb_resp_entry;
  reg [31:0] GEN_356;
  reg  ex_reg_btb_resp_bht_history;
  reg [31:0] GEN_357;
  reg [1:0] ex_reg_btb_resp_bht_value;
  reg [31:0] GEN_358;
  reg  ex_reg_xcpt;
  reg [31:0] GEN_359;
  reg  ex_reg_flush_pipe;
  reg [31:0] GEN_360;
  reg  ex_reg_load_use;
  reg [31:0] GEN_361;
  reg [31:0] ex_reg_cause;
  reg [31:0] GEN_362;
  reg  ex_reg_replay;
  reg [31:0] GEN_363;
  reg [31:0] ex_reg_pc;
  reg [31:0] GEN_364;
  reg [31:0] ex_reg_inst;
  reg [31:0] GEN_365;
  reg  mem_reg_xcpt_interrupt;
  reg [31:0] GEN_366;
  reg  mem_reg_valid;
  reg [31:0] GEN_367;
  reg  mem_reg_btb_hit;
  reg [31:0] GEN_368;
  reg  mem_reg_btb_resp_taken;
  reg [31:0] GEN_369;
  reg  mem_reg_btb_resp_mask;
  reg [31:0] GEN_370;
  reg  mem_reg_btb_resp_bridx;
  reg [31:0] GEN_371;
  reg [31:0] mem_reg_btb_resp_target;
  reg [31:0] GEN_372;
  reg  mem_reg_btb_resp_entry;
  reg [31:0] GEN_373;
  reg  mem_reg_btb_resp_bht_history;
  reg [31:0] GEN_374;
  reg [1:0] mem_reg_btb_resp_bht_value;
  reg [31:0] GEN_375;
  reg  mem_reg_xcpt;
  reg [31:0] GEN_376;
  reg  mem_reg_replay;
  reg [31:0] GEN_377;
  reg  mem_reg_flush_pipe;
  reg [31:0] GEN_378;
  reg [31:0] mem_reg_cause;
  reg [31:0] GEN_379;
  reg  mem_reg_slow_bypass;
  reg [31:0] GEN_380;
  reg  mem_reg_load;
  reg [31:0] GEN_381;
  reg  mem_reg_store;
  reg [31:0] GEN_382;
  reg [31:0] mem_reg_pc;
  reg [31:0] GEN_383;
  reg [31:0] mem_reg_inst;
  reg [31:0] GEN_384;
  reg [31:0] mem_reg_wdata;
  reg [31:0] GEN_385;
  reg [31:0] mem_reg_rs2;
  reg [31:0] GEN_386;
  wire  take_pc_mem;
  reg  wb_reg_valid;
  reg [31:0] GEN_387;
  reg  wb_reg_xcpt;
  reg [31:0] GEN_388;
  reg  wb_reg_mem_xcpt;
  reg [31:0] GEN_389;
  reg  wb_reg_replay;
  reg [31:0] GEN_390;
  reg [31:0] wb_reg_cause;
  reg [31:0] GEN_391;
  reg [31:0] wb_reg_pc;
  reg [31:0] GEN_392;
  reg [31:0] wb_reg_inst;
  reg [31:0] GEN_393;
  reg [31:0] wb_reg_wdata;
  reg [31:0] GEN_394;
  reg [31:0] wb_reg_rs2;
  reg [31:0] GEN_395;
  wire  take_pc_wb;
  wire  take_pc_mem_wb;
  wire  id_ctrl_legal;
  wire  id_ctrl_fp;
  wire  id_ctrl_rocc;
  wire  id_ctrl_branch;
  wire  id_ctrl_jal;
  wire  id_ctrl_jalr;
  wire  id_ctrl_rxs2;
  wire  id_ctrl_rxs1;
  wire [1:0] id_ctrl_sel_alu2;
  wire [1:0] id_ctrl_sel_alu1;
  wire [2:0] id_ctrl_sel_imm;
  wire  id_ctrl_alu_dw;
  wire [3:0] id_ctrl_alu_fn;
  wire  id_ctrl_mem;
  wire [4:0] id_ctrl_mem_cmd;
  wire [2:0] id_ctrl_mem_type;
  wire  id_ctrl_rfs1;
  wire  id_ctrl_rfs2;
  wire  id_ctrl_rfs3;
  wire  id_ctrl_wfd;
  wire  id_ctrl_div;
  wire  id_ctrl_wxd;
  wire [2:0] id_ctrl_csr;
  wire  id_ctrl_fence_i;
  wire  id_ctrl_fence;
  wire  id_ctrl_amo;
  wire [31:0] T_6562;
  wire  T_6564;
  wire [31:0] T_6566;
  wire  T_6568;
  wire [31:0] T_6570;
  wire  T_6572;
  wire [31:0] T_6574;
  wire  T_6576;
  wire [31:0] T_6578;
  wire  T_6580;
  wire [31:0] T_6582;
  wire  T_6584;
  wire [31:0] T_6586;
  wire  T_6588;
  wire [31:0] T_6590;
  wire  T_6592;
  wire [31:0] T_6594;
  wire  T_6596;
  wire [31:0] T_6598;
  wire  T_6600;
  wire  T_6604;
  wire  T_6608;
  wire [31:0] T_6610;
  wire  T_6612;
  wire  T_6616;
  wire  T_6618;
  wire  T_6620;
  wire  T_6622;
  wire [31:0] T_6624;
  wire  T_6626;
  wire [31:0] T_6628;
  wire  T_6630;
  wire [31:0] T_6632;
  wire  T_6634;
  wire  T_6638;
  wire  T_6641;
  wire  T_6642;
  wire  T_6643;
  wire  T_6644;
  wire  T_6645;
  wire  T_6646;
  wire  T_6647;
  wire  T_6648;
  wire  T_6649;
  wire  T_6650;
  wire  T_6651;
  wire  T_6652;
  wire  T_6653;
  wire  T_6654;
  wire  T_6655;
  wire  T_6656;
  wire  T_6657;
  wire  T_6658;
  wire  T_6659;
  wire  T_6660;
  wire [31:0] T_6664;
  wire  T_6666;
  wire [31:0] T_6670;
  wire  T_6672;
  wire [31:0] T_6676;
  wire  T_6678;
  wire [31:0] T_6682;
  wire  T_6684;
  wire [31:0] T_6686;
  wire  T_6688;
  wire  T_6691;
  wire [31:0] T_6693;
  wire  T_6695;
  wire [31:0] T_6697;
  wire  T_6699;
  wire [31:0] T_6701;
  wire  T_6703;
  wire  T_6706;
  wire  T_6707;
  wire [31:0] T_6709;
  wire  T_6711;
  wire [31:0] T_6713;
  wire  T_6715;
  wire [31:0] T_6717;
  wire  T_6719;
  wire [31:0] T_6721;
  wire  T_6723;
  wire  T_6726;
  wire  T_6727;
  wire  T_6728;
  wire [31:0] T_6730;
  wire  T_6732;
  wire [31:0] T_6734;
  wire  T_6736;
  wire  T_6739;
  wire  T_6740;
  wire [1:0] T_6741;
  wire [31:0] T_6747;
  wire  T_6749;
  wire [31:0] T_6751;
  wire  T_6753;
  wire  T_6756;
  wire [1:0] T_6757;
  wire  T_6761;
  wire  T_6764;
  wire  T_6768;
  wire  T_6771;
  wire  T_6775;
  wire [31:0] T_6777;
  wire  T_6779;
  wire  T_6782;
  wire  T_6783;
  wire [1:0] T_6784;
  wire [2:0] T_6785;
  wire [31:0] T_6793;
  wire  T_6795;
  wire [31:0] T_6797;
  wire  T_6799;
  wire [31:0] T_6801;
  wire  T_6803;
  wire  T_6806;
  wire  T_6807;
  wire [31:0] T_6809;
  wire  T_6811;
  wire [31:0] T_6813;
  wire  T_6815;
  wire [31:0] T_6817;
  wire  T_6819;
  wire [31:0] T_6821;
  wire  T_6823;
  wire [31:0] T_6825;
  wire  T_6827;
  wire [31:0] T_6829;
  wire  T_6831;
  wire  T_6834;
  wire  T_6835;
  wire  T_6836;
  wire  T_6837;
  wire  T_6838;
  wire [31:0] T_6840;
  wire  T_6842;
  wire [31:0] T_6844;
  wire  T_6846;
  wire [31:0] T_6848;
  wire  T_6850;
  wire [31:0] T_6852;
  wire  T_6854;
  wire  T_6857;
  wire  T_6858;
  wire  T_6859;
  wire [31:0] T_6861;
  wire  T_6863;
  wire [31:0] T_6865;
  wire  T_6867;
  wire  T_6870;
  wire  T_6871;
  wire  T_6872;
  wire [1:0] T_6873;
  wire [2:0] T_6874;
  wire [3:0] T_6875;
  wire [31:0] T_6877;
  wire  T_6879;
  wire [31:0] T_6881;
  wire  T_6883;
  wire  T_6886;
  wire  T_6887;
  wire  T_6888;
  wire  T_6892;
  wire  T_6895;
  wire [1:0] T_6901;
  wire [2:0] T_6902;
  wire [3:0] T_6903;
  wire [4:0] T_6904;
  wire [31:0] T_6906;
  wire  T_6908;
  wire [31:0] T_6912;
  wire  T_6914;
  wire [31:0] T_6918;
  wire  T_6920;
  wire [1:0] T_6923;
  wire [2:0] T_6924;
  wire [31:0] T_6930;
  wire  T_6932;
  wire [31:0] T_6936;
  wire  T_6938;
  wire [31:0] T_6940;
  wire  T_6942;
  wire  T_6946;
  wire [31:0] T_6948;
  wire  T_6950;
  wire [31:0] T_6952;
  wire  T_6954;
  wire  T_6957;
  wire  T_6958;
  wire  T_6959;
  wire  T_6960;
  wire  T_6961;
  wire [31:0] T_6963;
  wire  T_6965;
  wire [31:0] T_6969;
  wire  T_6971;
  wire [31:0] T_6975;
  wire  T_6977;
  wire [1:0] T_6980;
  wire [2:0] T_6981;
  wire [31:0] T_6983;
  wire  T_6985;
  wire  T_6991;
  wire [4:0] id_raddr3;
  wire [4:0] id_raddr2;
  wire [4:0] id_raddr1;
  wire [4:0] id_waddr;
  wire  id_load_use;
  reg  id_reg_fence;
  reg [31:0] GEN_396;
  reg [31:0] T_6999 [0:30];
  reg [31:0] GEN_397;
  wire [31:0] T_6999_T_7009_data;
  wire [4:0] T_6999_T_7009_addr;
  wire  T_6999_T_7009_en;
  reg [31:0] GEN_398;
  wire [31:0] T_6999_T_7020_data;
  wire [4:0] T_6999_T_7020_addr;
  wire  T_6999_T_7020_en;
  reg [31:0] GEN_399;
  wire [31:0] T_6999_T_7648_data;
  wire [4:0] T_6999_T_7648_addr;
  wire  T_6999_T_7648_mask;
  wire  T_6999_T_7648_en;
  wire [31:0] T_7001;
  wire  T_7004;
  wire [4:0] T_7008;
  wire [31:0] T_7010;
  wire [31:0] T_7012;
  wire [4:0] T_7019;
  wire [31:0] T_7021;
  wire  ctrl_killd;
  wire  csr_clk;
  wire  csr_reset;
  wire  csr_io_prci_reset;
  wire  csr_io_prci_id;
  wire  csr_io_prci_interrupts_meip;
  wire  csr_io_prci_interrupts_seip;
  wire  csr_io_prci_interrupts_debug;
  wire  csr_io_prci_interrupts_mtip;
  wire  csr_io_prci_interrupts_msip;
  wire [11:0] csr_io_rw_addr;
  wire [2:0] csr_io_rw_cmd;
  wire [31:0] csr_io_rw_rdata;
  wire [31:0] csr_io_rw_wdata;
  wire  csr_io_csr_stall;
  wire  csr_io_csr_xcpt;
  wire  csr_io_eret;
  wire  csr_io_singleStep;
  wire  csr_io_status_debug;
  wire [1:0] csr_io_status_prv;
  wire  csr_io_status_sd;
  wire [30:0] csr_io_status_zero3;
  wire  csr_io_status_sd_rv32;
  wire [1:0] csr_io_status_zero2;
  wire [4:0] csr_io_status_vm;
  wire [3:0] csr_io_status_zero1;
  wire  csr_io_status_mxr;
  wire  csr_io_status_pum;
  wire  csr_io_status_mprv;
  wire [1:0] csr_io_status_xs;
  wire [1:0] csr_io_status_fs;
  wire [1:0] csr_io_status_mpp;
  wire [1:0] csr_io_status_hpp;
  wire  csr_io_status_spp;
  wire  csr_io_status_mpie;
  wire  csr_io_status_hpie;
  wire  csr_io_status_spie;
  wire  csr_io_status_upie;
  wire  csr_io_status_mie;
  wire  csr_io_status_hie;
  wire  csr_io_status_sie;
  wire  csr_io_status_uie;
  wire [6:0] csr_io_ptbr_asid;
  wire [21:0] csr_io_ptbr_ppn;
  wire [31:0] csr_io_evec;
  wire  csr_io_exception;
  wire  csr_io_retire;
  wire [31:0] csr_io_cause;
  wire [31:0] csr_io_pc;
  wire [31:0] csr_io_badaddr;
  wire  csr_io_fatc;
  wire [31:0] csr_io_time;
  wire [2:0] csr_io_fcsr_rm;
  wire  csr_io_fcsr_flags_valid;
  wire [4:0] csr_io_fcsr_flags_bits;
  wire  csr_io_rocc_cmd_ready;
  wire  csr_io_rocc_cmd_valid;
  wire [6:0] csr_io_rocc_cmd_bits_inst_funct;
  wire [4:0] csr_io_rocc_cmd_bits_inst_rs2;
  wire [4:0] csr_io_rocc_cmd_bits_inst_rs1;
  wire  csr_io_rocc_cmd_bits_inst_xd;
  wire  csr_io_rocc_cmd_bits_inst_xs1;
  wire  csr_io_rocc_cmd_bits_inst_xs2;
  wire [4:0] csr_io_rocc_cmd_bits_inst_rd;
  wire [6:0] csr_io_rocc_cmd_bits_inst_opcode;
  wire [31:0] csr_io_rocc_cmd_bits_rs1;
  wire [31:0] csr_io_rocc_cmd_bits_rs2;
  wire  csr_io_rocc_cmd_bits_status_debug;
  wire [1:0] csr_io_rocc_cmd_bits_status_prv;
  wire  csr_io_rocc_cmd_bits_status_sd;
  wire [30:0] csr_io_rocc_cmd_bits_status_zero3;
  wire  csr_io_rocc_cmd_bits_status_sd_rv32;
  wire [1:0] csr_io_rocc_cmd_bits_status_zero2;
  wire [4:0] csr_io_rocc_cmd_bits_status_vm;
  wire [3:0] csr_io_rocc_cmd_bits_status_zero1;
  wire  csr_io_rocc_cmd_bits_status_mxr;
  wire  csr_io_rocc_cmd_bits_status_pum;
  wire  csr_io_rocc_cmd_bits_status_mprv;
  wire [1:0] csr_io_rocc_cmd_bits_status_xs;
  wire [1:0] csr_io_rocc_cmd_bits_status_fs;
  wire [1:0] csr_io_rocc_cmd_bits_status_mpp;
  wire [1:0] csr_io_rocc_cmd_bits_status_hpp;
  wire  csr_io_rocc_cmd_bits_status_spp;
  wire  csr_io_rocc_cmd_bits_status_mpie;
  wire  csr_io_rocc_cmd_bits_status_hpie;
  wire  csr_io_rocc_cmd_bits_status_spie;
  wire  csr_io_rocc_cmd_bits_status_upie;
  wire  csr_io_rocc_cmd_bits_status_mie;
  wire  csr_io_rocc_cmd_bits_status_hie;
  wire  csr_io_rocc_cmd_bits_status_sie;
  wire  csr_io_rocc_cmd_bits_status_uie;
  wire  csr_io_rocc_resp_ready;
  wire  csr_io_rocc_resp_valid;
  wire [4:0] csr_io_rocc_resp_bits_rd;
  wire [31:0] csr_io_rocc_resp_bits_data;
  wire  csr_io_rocc_mem_req_ready;
  wire  csr_io_rocc_mem_req_valid;
  wire [31:0] csr_io_rocc_mem_req_bits_addr;
  wire [8:0] csr_io_rocc_mem_req_bits_tag;
  wire [4:0] csr_io_rocc_mem_req_bits_cmd;
  wire [2:0] csr_io_rocc_mem_req_bits_typ;
  wire  csr_io_rocc_mem_req_bits_phys;
  wire [31:0] csr_io_rocc_mem_req_bits_data;
  wire  csr_io_rocc_mem_s1_kill;
  wire [31:0] csr_io_rocc_mem_s1_data;
  wire  csr_io_rocc_mem_s2_nack;
  wire  csr_io_rocc_mem_resp_valid;
  wire [31:0] csr_io_rocc_mem_resp_bits_addr;
  wire [8:0] csr_io_rocc_mem_resp_bits_tag;
  wire [4:0] csr_io_rocc_mem_resp_bits_cmd;
  wire [2:0] csr_io_rocc_mem_resp_bits_typ;
  wire [31:0] csr_io_rocc_mem_resp_bits_data;
  wire  csr_io_rocc_mem_resp_bits_replay;
  wire  csr_io_rocc_mem_resp_bits_has_data;
  wire [31:0] csr_io_rocc_mem_resp_bits_data_word_bypass;
  wire [31:0] csr_io_rocc_mem_resp_bits_store_data;
  wire  csr_io_rocc_mem_replay_next;
  wire  csr_io_rocc_mem_xcpt_ma_ld;
  wire  csr_io_rocc_mem_xcpt_ma_st;
  wire  csr_io_rocc_mem_xcpt_pf_ld;
  wire  csr_io_rocc_mem_xcpt_pf_st;
  wire  csr_io_rocc_mem_invalidate_lr;
  wire  csr_io_rocc_mem_ordered;
  wire  csr_io_rocc_busy;
  wire  csr_io_rocc_interrupt;
  wire  csr_io_rocc_autl_acquire_ready;
  wire  csr_io_rocc_autl_acquire_valid;
  wire [25:0] csr_io_rocc_autl_acquire_bits_addr_block;
  wire  csr_io_rocc_autl_acquire_bits_client_xact_id;
  wire [2:0] csr_io_rocc_autl_acquire_bits_addr_beat;
  wire  csr_io_rocc_autl_acquire_bits_is_builtin_type;
  wire [2:0] csr_io_rocc_autl_acquire_bits_a_type;
  wire [11:0] csr_io_rocc_autl_acquire_bits_union;
  wire [63:0] csr_io_rocc_autl_acquire_bits_data;
  wire  csr_io_rocc_autl_grant_ready;
  wire  csr_io_rocc_autl_grant_valid;
  wire [2:0] csr_io_rocc_autl_grant_bits_addr_beat;
  wire  csr_io_rocc_autl_grant_bits_client_xact_id;
  wire [1:0] csr_io_rocc_autl_grant_bits_manager_xact_id;
  wire  csr_io_rocc_autl_grant_bits_is_builtin_type;
  wire [3:0] csr_io_rocc_autl_grant_bits_g_type;
  wire [63:0] csr_io_rocc_autl_grant_bits_data;
  wire  csr_io_rocc_fpu_req_ready;
  wire  csr_io_rocc_fpu_req_valid;
  wire [4:0] csr_io_rocc_fpu_req_bits_cmd;
  wire  csr_io_rocc_fpu_req_bits_ldst;
  wire  csr_io_rocc_fpu_req_bits_wen;
  wire  csr_io_rocc_fpu_req_bits_ren1;
  wire  csr_io_rocc_fpu_req_bits_ren2;
  wire  csr_io_rocc_fpu_req_bits_ren3;
  wire  csr_io_rocc_fpu_req_bits_swap12;
  wire  csr_io_rocc_fpu_req_bits_swap23;
  wire  csr_io_rocc_fpu_req_bits_single;
  wire  csr_io_rocc_fpu_req_bits_fromint;
  wire  csr_io_rocc_fpu_req_bits_toint;
  wire  csr_io_rocc_fpu_req_bits_fastpipe;
  wire  csr_io_rocc_fpu_req_bits_fma;
  wire  csr_io_rocc_fpu_req_bits_div;
  wire  csr_io_rocc_fpu_req_bits_sqrt;
  wire  csr_io_rocc_fpu_req_bits_round;
  wire  csr_io_rocc_fpu_req_bits_wflags;
  wire [2:0] csr_io_rocc_fpu_req_bits_rm;
  wire [1:0] csr_io_rocc_fpu_req_bits_typ;
  wire [64:0] csr_io_rocc_fpu_req_bits_in1;
  wire [64:0] csr_io_rocc_fpu_req_bits_in2;
  wire [64:0] csr_io_rocc_fpu_req_bits_in3;
  wire  csr_io_rocc_fpu_resp_ready;
  wire  csr_io_rocc_fpu_resp_valid;
  wire [64:0] csr_io_rocc_fpu_resp_bits_data;
  wire [4:0] csr_io_rocc_fpu_resp_bits_exc;
  wire  csr_io_rocc_exception;
  wire [11:0] csr_io_rocc_csr_waddr;
  wire [31:0] csr_io_rocc_csr_wdata;
  wire  csr_io_rocc_csr_wen;
  wire  csr_io_rocc_host_id;
  wire  csr_io_interrupt;
  wire [31:0] csr_io_interrupt_cause;
  wire [3:0] csr_io_bp_0_control_tdrtype;
  wire [4:0] csr_io_bp_0_control_bpamaskmax;
  wire [3:0] csr_io_bp_0_control_reserved;
  wire [7:0] csr_io_bp_0_control_bpaction;
  wire [3:0] csr_io_bp_0_control_bpmatch;
  wire  csr_io_bp_0_control_m;
  wire  csr_io_bp_0_control_h;
  wire  csr_io_bp_0_control_s;
  wire  csr_io_bp_0_control_u;
  wire  csr_io_bp_0_control_r;
  wire  csr_io_bp_0_control_w;
  wire  csr_io_bp_0_control_x;
  wire [31:0] csr_io_bp_0_address;
  wire [3:0] csr_io_bp_1_control_tdrtype;
  wire [4:0] csr_io_bp_1_control_bpamaskmax;
  wire [3:0] csr_io_bp_1_control_reserved;
  wire [7:0] csr_io_bp_1_control_bpaction;
  wire [3:0] csr_io_bp_1_control_bpmatch;
  wire  csr_io_bp_1_control_m;
  wire  csr_io_bp_1_control_h;
  wire  csr_io_bp_1_control_s;
  wire  csr_io_bp_1_control_u;
  wire  csr_io_bp_1_control_r;
  wire  csr_io_bp_1_control_w;
  wire  csr_io_bp_1_control_x;
  wire [31:0] csr_io_bp_1_address;
  wire  id_csr_en;
  wire  id_system_insn;
  wire  T_7023;
  wire  T_7024;
  wire  T_7025;
  wire  id_csr_ren;
  wire [2:0] id_csr;
  wire [11:0] id_csr_addr;
  wire  T_7029;
  wire  T_7030;
  wire [11:0] T_7084;
  wire  T_7086;
  wire [11:0] T_7088;
  wire  T_7090;
  wire  T_7093;
  wire  T_7096;
  wire  T_7097;
  wire  id_csr_flush;
  wire  T_7099;
  wire  T_7101;
  wire  T_7103;
  wire  T_7104;
  wire  T_7105;
  wire  T_7107;
  wire  T_7109;
  wire  T_7110;
  wire  id_illegal_insn;
  wire  id_amo_aq;
  wire  id_amo_rl;
  wire  T_7111;
  wire  id_fence_next;
  wire  T_7113;
  wire  id_mem_busy;
  wire  T_7119;
  wire  T_7121;
  wire  T_7122;
  wire  T_7124;
  wire  T_7125;
  wire  T_7126;
  wire  T_7127;
  wire  T_7128;
  wire  T_7129;
  wire  T_7130;
  wire  bpu_clk;
  wire  bpu_reset;
  wire  bpu_io_status_debug;
  wire [1:0] bpu_io_status_prv;
  wire  bpu_io_status_sd;
  wire [30:0] bpu_io_status_zero3;
  wire  bpu_io_status_sd_rv32;
  wire [1:0] bpu_io_status_zero2;
  wire [4:0] bpu_io_status_vm;
  wire [3:0] bpu_io_status_zero1;
  wire  bpu_io_status_mxr;
  wire  bpu_io_status_pum;
  wire  bpu_io_status_mprv;
  wire [1:0] bpu_io_status_xs;
  wire [1:0] bpu_io_status_fs;
  wire [1:0] bpu_io_status_mpp;
  wire [1:0] bpu_io_status_hpp;
  wire  bpu_io_status_spp;
  wire  bpu_io_status_mpie;
  wire  bpu_io_status_hpie;
  wire  bpu_io_status_spie;
  wire  bpu_io_status_upie;
  wire  bpu_io_status_mie;
  wire  bpu_io_status_hie;
  wire  bpu_io_status_sie;
  wire  bpu_io_status_uie;
  wire [3:0] bpu_io_bp_0_control_tdrtype;
  wire [4:0] bpu_io_bp_0_control_bpamaskmax;
  wire [3:0] bpu_io_bp_0_control_reserved;
  wire [7:0] bpu_io_bp_0_control_bpaction;
  wire [3:0] bpu_io_bp_0_control_bpmatch;
  wire  bpu_io_bp_0_control_m;
  wire  bpu_io_bp_0_control_h;
  wire  bpu_io_bp_0_control_s;
  wire  bpu_io_bp_0_control_u;
  wire  bpu_io_bp_0_control_r;
  wire  bpu_io_bp_0_control_w;
  wire  bpu_io_bp_0_control_x;
  wire [31:0] bpu_io_bp_0_address;
  wire [3:0] bpu_io_bp_1_control_tdrtype;
  wire [4:0] bpu_io_bp_1_control_bpamaskmax;
  wire [3:0] bpu_io_bp_1_control_reserved;
  wire [7:0] bpu_io_bp_1_control_bpaction;
  wire [3:0] bpu_io_bp_1_control_bpmatch;
  wire  bpu_io_bp_1_control_m;
  wire  bpu_io_bp_1_control_h;
  wire  bpu_io_bp_1_control_s;
  wire  bpu_io_bp_1_control_u;
  wire  bpu_io_bp_1_control_r;
  wire  bpu_io_bp_1_control_w;
  wire  bpu_io_bp_1_control_x;
  wire [31:0] bpu_io_bp_1_address;
  wire [31:0] bpu_io_pc;
  wire [31:0] bpu_io_ea;
  wire  bpu_io_xcpt_if;
  wire  bpu_io_xcpt_ld;
  wire  bpu_io_xcpt_st;
  wire  T_7134;
  wire  T_7135;
  wire  id_xcpt;
  wire [1:0] T_7136;
  wire [1:0] T_7137;
  wire [31:0] id_cause;
  wire [4:0] ex_waddr;
  wire [4:0] mem_waddr;
  wire [4:0] wb_waddr;
  wire  T_7141;
  wire  T_7142;
  wire  T_7144;
  wire  T_7145;
  wire  T_7147;
  wire  T_7149;
  wire  T_7150;
  wire  T_7151;
  wire  T_7152;
  wire  T_7154;
  wire  T_7155;
  wire  T_7157;
  wire  T_7158;
  wire  T_7159;
  wire  T_7160;
  wire  T_7162;
  wire [31:0] bypass_mux_0;
  wire [31:0] bypass_mux_1;
  wire [31:0] bypass_mux_2;
  wire [31:0] bypass_mux_3;
  reg  ex_reg_rs_bypass_0;
  reg [31:0] GEN_400;
  reg  ex_reg_rs_bypass_1;
  reg [31:0] GEN_401;
  reg [1:0] ex_reg_rs_lsb_0;
  reg [31:0] GEN_402;
  reg [1:0] ex_reg_rs_lsb_1;
  reg [31:0] GEN_403;
  reg [29:0] ex_reg_rs_msb_0;
  reg [31:0] GEN_404;
  reg [29:0] ex_reg_rs_msb_1;
  reg [31:0] GEN_405;
  wire [31:0] T_7190;
  wire [31:0] GEN_0;
  wire [31:0] GEN_2;
  wire [31:0] GEN_3;
  wire [31:0] GEN_4;
  wire [31:0] T_7191;
  wire [31:0] T_7192;
  wire [31:0] GEN_1;
  wire [31:0] GEN_5;
  wire [31:0] GEN_6;
  wire [31:0] GEN_7;
  wire [31:0] T_7193;
  wire  T_7194;
  wire  T_7196;
  wire  T_7197;
  wire  T_7198;
  wire  T_7199;
  wire [10:0] T_7200;
  wire [10:0] T_7201;
  wire [10:0] T_7202;
  wire  T_7203;
  wire  T_7204;
  wire  T_7205;
  wire [7:0] T_7206;
  wire [7:0] T_7207;
  wire [7:0] T_7208;
  wire  T_7211;
  wire  T_7213;
  wire  T_7214;
  wire  T_7215;
  wire  T_7216;
  wire  T_7217;
  wire  T_7218;
  wire  T_7219;
  wire  T_7220;
  wire  T_7221;
  wire [5:0] T_7226;
  wire [5:0] T_7227;
  wire  T_7230;
  wire  T_7232;
  wire [3:0] T_7233;
  wire [3:0] T_7235;
  wire [3:0] T_7236;
  wire [3:0] T_7237;
  wire [3:0] T_7238;
  wire [3:0] T_7239;
  wire  T_7242;
  wire  T_7245;
  wire  T_7248;
  wire  T_7250;
  wire  T_7252;
  wire [9:0] T_7253;
  wire [10:0] T_7254;
  wire  T_7255;
  wire [7:0] T_7256;
  wire [8:0] T_7257;
  wire [10:0] T_7258;
  wire  T_7259;
  wire [11:0] T_7260;
  wire [20:0] T_7261;
  wire [31:0] T_7262;
  wire [31:0] ex_imm;
  wire [31:0] T_7264;
  wire [31:0] T_7265;
  wire  T_7266;
  wire [31:0] T_7267;
  wire  T_7268;
  wire [31:0] ex_op1;
  wire [31:0] T_7270;
  wire  T_7272;
  wire [3:0] T_7273;
  wire  T_7274;
  wire [31:0] T_7275;
  wire  T_7276;
  wire [31:0] ex_op2;
  wire  alu_clk;
  wire  alu_reset;
  wire  alu_io_dw;
  wire [3:0] alu_io_fn;
  wire [31:0] alu_io_in2;
  wire [31:0] alu_io_in1;
  wire [31:0] alu_io_out;
  wire [31:0] alu_io_adder_out;
  wire  alu_io_cmp_out;
  wire [31:0] T_7277;
  wire [31:0] T_7278;
  wire  div_clk;
  wire  div_reset;
  wire  div_io_req_ready;
  wire  div_io_req_valid;
  wire [3:0] div_io_req_bits_fn;
  wire  div_io_req_bits_dw;
  wire [31:0] div_io_req_bits_in1;
  wire [31:0] div_io_req_bits_in2;
  wire [4:0] div_io_req_bits_tag;
  wire  div_io_kill;
  wire  div_io_resp_ready;
  wire  div_io_resp_valid;
  wire [31:0] div_io_resp_bits_data;
  wire [4:0] div_io_resp_bits_tag;
  wire  T_7279;
  wire  T_7281;
  wire  T_7283;
  wire  T_7284;
  wire  T_7285;
  wire  T_7288;
  wire  T_7292;
  wire [31:0] GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire [31:0] GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire [1:0] GEN_15;
  wire  T_7295;
  wire  T_7296;
  wire  T_7297;
  wire  GEN_16;
  wire  GEN_17;
  wire  T_7300;
  wire  T_7301;
  wire  T_7302;
  wire [1:0] T_7307;
  wire [1:0] T_7308;
  wire [1:0] T_7309;
  wire  T_7311;
  wire  T_7312;
  wire [1:0] T_7313;
  wire [29:0] T_7314;
  wire [1:0] GEN_18;
  wire [29:0] GEN_19;
  wire  T_7315;
  wire  T_7316;
  wire  T_7317;
  wire [1:0] T_7322;
  wire [1:0] T_7323;
  wire [1:0] T_7324;
  wire  T_7326;
  wire  T_7327;
  wire [1:0] T_7328;
  wire [29:0] T_7329;
  wire [1:0] GEN_20;
  wire [29:0] GEN_21;
  wire  GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_29;
  wire [1:0] GEN_30;
  wire [1:0] GEN_31;
  wire [2:0] GEN_32;
  wire  GEN_33;
  wire [3:0] GEN_34;
  wire  GEN_35;
  wire [4:0] GEN_36;
  wire [2:0] GEN_37;
  wire  GEN_38;
  wire  GEN_39;
  wire  GEN_40;
  wire  GEN_41;
  wire  GEN_42;
  wire  GEN_43;
  wire [2:0] GEN_44;
  wire  GEN_45;
  wire  GEN_46;
  wire  GEN_47;
  wire  GEN_48;
  wire  GEN_49;
  wire  GEN_50;
  wire  GEN_51;
  wire [31:0] GEN_52;
  wire  GEN_53;
  wire  GEN_54;
  wire [1:0] GEN_55;
  wire  GEN_56;
  wire  GEN_57;
  wire  GEN_58;
  wire [1:0] GEN_59;
  wire [29:0] GEN_60;
  wire  GEN_61;
  wire [1:0] GEN_62;
  wire [29:0] GEN_63;
  wire  T_7332;
  wire  T_7333;
  wire [31:0] GEN_64;
  wire [31:0] GEN_65;
  wire  T_7334;
  wire  ex_pc_valid;
  wire  T_7336;
  wire  wb_dcache_miss;
  wire  T_7338;
  wire  T_7339;
  wire  T_7341;
  wire  T_7342;
  wire  replay_ex_structural;
  wire  replay_ex_load_use;
  wire  T_7343;
  wire  T_7344;
  wire  replay_ex;
  wire  T_7345;
  wire  T_7347;
  wire  ctrl_killx;
  wire  T_7348;
  wire [2:0] T_7354_0;
  wire [2:0] T_7354_1;
  wire [2:0] T_7354_2;
  wire [2:0] T_7354_3;
  wire  T_7356;
  wire  T_7357;
  wire  T_7358;
  wire  T_7359;
  wire  T_7362;
  wire  T_7363;
  wire  T_7364;
  wire  ex_slow_bypass;
  wire  T_7365;
  wire  T_7366;
  wire  ex_xcpt;
  wire [31:0] ex_cause;
  wire  mem_br_taken;
  wire [31:0] T_7368;
  wire  T_7369;
  wire  T_7372;
  wire  T_7373;
  wire [10:0] T_7378;
  wire [7:0] T_7382;
  wire [7:0] T_7383;
  wire [7:0] T_7384;
  wire  T_7390;
  wire  T_7391;
  wire  T_7393;
  wire  T_7394;
  wire [5:0] T_7402;
  wire [3:0] T_7409;
  wire [3:0] T_7412;
  wire [9:0] T_7429;
  wire [10:0] T_7430;
  wire  T_7431;
  wire [7:0] T_7432;
  wire [8:0] T_7433;
  wire [10:0] T_7434;
  wire  T_7435;
  wire [11:0] T_7436;
  wire [20:0] T_7437;
  wire [31:0] T_7438;
  wire [31:0] T_7439;
  wire [9:0] T_7499;
  wire [10:0] T_7500;
  wire  T_7501;
  wire [7:0] T_7502;
  wire [8:0] T_7503;
  wire [20:0] T_7507;
  wire [31:0] T_7508;
  wire [31:0] T_7509;
  wire [31:0] T_7511;
  wire [31:0] T_7512;
  wire [32:0] T_7513;
  wire [31:0] T_7514;
  wire [31:0] mem_br_target;
  wire [31:0] T_7515;
  wire [31:0] T_7516;
  wire [31:0] mem_int_wdata;
  wire [31:0] T_7518;
  wire [31:0] T_7520;
  wire [31:0] T_7521;
  wire [31:0] mem_npc;
  wire  T_7522;
  wire  T_7523;
  wire  T_7525;
  wire  mem_wrong_npc;
  wire  mem_npc_misaligned;
  wire  T_7528;
  wire  mem_misprediction;
  wire  T_7529;
  wire  want_take_pc_mem;
  wire  T_7531;
  wire  T_7532;
  wire  T_7534;
  wire  T_7537;
  wire  T_7540;
  wire  T_7543;
  wire [31:0] GEN_66;
  wire  T_7544;
  wire  T_7545;
  wire  T_7546;
  wire  T_7548;
  wire  T_7549;
  wire  T_7550;
  wire  T_7551;
  wire  T_7552;
  wire  T_7553;
  wire  T_7554;
  wire  T_7556;
  wire  T_7560;
  wire  T_7561;
  wire  GEN_67;
  wire  GEN_68;
  wire  GEN_69;
  wire [31:0] GEN_70;
  wire  GEN_71;
  wire  GEN_72;
  wire [1:0] GEN_73;
  wire  T_7562;
  wire  T_7563;
  wire [31:0] GEN_74;
  wire  GEN_75;
  wire  GEN_76;
  wire  GEN_77;
  wire  GEN_78;
  wire  GEN_79;
  wire  GEN_80;
  wire  GEN_81;
  wire  GEN_82;
  wire [1:0] GEN_83;
  wire [1:0] GEN_84;
  wire [2:0] GEN_85;
  wire  GEN_86;
  wire [3:0] GEN_87;
  wire  GEN_88;
  wire [4:0] GEN_89;
  wire [2:0] GEN_90;
  wire  GEN_91;
  wire  GEN_92;
  wire  GEN_93;
  wire  GEN_94;
  wire  GEN_95;
  wire  GEN_96;
  wire [2:0] GEN_97;
  wire  GEN_98;
  wire  GEN_99;
  wire  GEN_100;
  wire  GEN_101;
  wire  GEN_102;
  wire  GEN_103;
  wire  GEN_104;
  wire  GEN_105;
  wire  GEN_106;
  wire [31:0] GEN_107;
  wire  GEN_108;
  wire  GEN_109;
  wire [1:0] GEN_110;
  wire  GEN_111;
  wire  GEN_112;
  wire [31:0] GEN_113;
  wire [31:0] GEN_114;
  wire [31:0] GEN_115;
  wire [31:0] GEN_116;
  wire  T_7564;
  wire  T_7566;
  wire  T_7568;
  wire  T_7570;
  wire  T_7572;
  wire  T_7574;
  wire  T_7576;
  wire  T_7578;
  wire  T_7579;
  wire  T_7580;
  wire  T_7581;
  wire  T_7582;
  wire  mem_new_xcpt;
  wire [2:0] T_7583;
  wire [2:0] T_7584;
  wire [2:0] T_7585;
  wire [2:0] T_7586;
  wire [2:0] T_7587;
  wire [2:0] mem_new_cause;
  wire  T_7588;
  wire  T_7589;
  wire  mem_xcpt;
  wire [31:0] mem_cause;
  wire  dcache_kill_mem;
  wire  T_7591;
  wire  fpu_kill_mem;
  wire  T_7592;
  wire  replay_mem;
  wire  T_7593;
  wire  T_7594;
  wire  T_7596;
  wire  killm_common;
  wire  T_7597;
  reg  T_7598;
  reg [31:0] GEN_406;
  wire  T_7599;
  wire  T_7600;
  wire  ctrl_killm;
  wire  T_7602;
  wire  T_7604;
  wire  T_7605;
  wire  T_7608;
  wire  T_7612;
  wire  T_7613;
  wire [31:0] GEN_117;
  wire  T_7614;
  wire  T_7615;
  wire  T_7616;
  wire [31:0] T_7617;
  wire [31:0] GEN_118;
  wire  GEN_119;
  wire  GEN_120;
  wire  GEN_121;
  wire  GEN_122;
  wire  GEN_123;
  wire  GEN_124;
  wire  GEN_125;
  wire  GEN_126;
  wire [1:0] GEN_127;
  wire [1:0] GEN_128;
  wire [2:0] GEN_129;
  wire  GEN_130;
  wire [3:0] GEN_131;
  wire  GEN_132;
  wire [4:0] GEN_133;
  wire [2:0] GEN_134;
  wire  GEN_135;
  wire  GEN_136;
  wire  GEN_137;
  wire  GEN_138;
  wire  GEN_139;
  wire  GEN_140;
  wire [2:0] GEN_141;
  wire  GEN_142;
  wire  GEN_143;
  wire  GEN_144;
  wire [31:0] GEN_145;
  wire [31:0] GEN_146;
  wire [31:0] GEN_147;
  wire [31:0] GEN_148;
  wire  T_7618;
  wire  wb_set_sboard;
  wire  replay_wb_common;
  wire  T_7621;
  wire  replay_wb_rocc;
  wire  replay_wb;
  wire  wb_xcpt;
  wire  T_7622;
  wire  T_7623;
  wire  T_7624;
  wire  dmem_resp_xpu;
  wire [7:0] dmem_resp_waddr;
  wire  dmem_resp_valid;
  wire  dmem_resp_replay;
  wire  T_7628;
  wire  T_7630;
  wire [31:0] ll_wdata;
  wire [7:0] ll_waddr;
  wire  T_7631;
  wire  ll_wen;
  wire  T_7632;
  wire  GEN_149;
  wire [7:0] GEN_150;
  wire  GEN_151;
  wire  T_7636;
  wire  T_7637;
  wire  T_7639;
  wire  wb_valid;
  wire  wb_wen;
  wire  rf_wen;
  wire [7:0] rf_waddr;
  wire  T_7640;
  wire  T_7641;
  wire [31:0] T_7642;
  wire [31:0] T_7643;
  wire [31:0] rf_wdata;
  wire  T_7645;
  wire [4:0] T_7646;
  wire [4:0] T_7647;
  wire [7:0] GEN_170;
  wire  T_7649;
  wire [31:0] GEN_152;
  wire [7:0] GEN_171;
  wire  T_7650;
  wire [31:0] GEN_153;
  wire [31:0] GEN_159;
  wire [31:0] GEN_160;
  wire  GEN_163;
  wire [31:0] GEN_166;
  wire [31:0] GEN_167;
  wire [31:0] T_7651;
  wire [11:0] T_7652;
  wire [2:0] T_7653;
  wire  T_7655;
  wire  T_7656;
  wire  T_7658;
  wire  T_7659;
  wire  T_7661;
  wire  T_7662;
  reg [31:0] T_7664;
  reg [31:0] GEN_407;
  wire [255:0] T_7667;
  wire [255:0] T_7669;
  wire [255:0] T_7670;
  wire [255:0] GEN_172;
  wire [255:0] T_7671;
  wire [255:0] GEN_168;
  wire [31:0] T_7673;
  wire  T_7674;
  wire  T_7675;
  wire [31:0] T_7676;
  wire  T_7677;
  wire  T_7678;
  wire [31:0] T_7679;
  wire  T_7680;
  wire  T_7681;
  wire  T_7682;
  wire  id_sboard_hazard;
  wire  T_7683;
  wire [31:0] T_7685;
  wire [31:0] T_7687;
  wire [255:0] GEN_173;
  wire [255:0] T_7688;
  wire  T_7689;
  wire [255:0] GEN_169;
  wire  T_7690;
  wire  T_7691;
  wire  T_7692;
  wire  T_7693;
  wire  T_7694;
  wire  ex_cannot_bypass;
  wire  T_7695;
  wire  T_7696;
  wire  T_7697;
  wire  T_7698;
  wire  T_7699;
  wire  T_7700;
  wire  T_7701;
  wire  T_7702;
  wire  data_hazard_ex;
  wire  T_7704;
  wire  T_7706;
  wire  T_7707;
  wire  T_7708;
  wire  T_7710;
  wire  T_7711;
  wire  T_7712;
  wire  T_7713;
  wire  fp_data_hazard_ex;
  wire  T_7714;
  wire  T_7715;
  wire  id_ex_hazard;
  wire  T_7717;
  wire  T_7718;
  wire  T_7719;
  wire  T_7720;
  wire  T_7721;
  wire  mem_cannot_bypass;
  wire  T_7722;
  wire  T_7723;
  wire  T_7724;
  wire  T_7725;
  wire  T_7726;
  wire  T_7727;
  wire  T_7728;
  wire  T_7729;
  wire  data_hazard_mem;
  wire  T_7731;
  wire  T_7733;
  wire  T_7734;
  wire  T_7735;
  wire  T_7737;
  wire  T_7738;
  wire  T_7739;
  wire  T_7740;
  wire  fp_data_hazard_mem;
  wire  T_7741;
  wire  T_7742;
  wire  id_mem_hazard;
  wire  T_7743;
  wire  T_7744;
  wire  T_7745;
  wire  T_7746;
  wire  T_7747;
  wire  T_7748;
  wire  T_7749;
  wire  T_7750;
  wire  T_7751;
  wire  T_7752;
  wire  data_hazard_wb;
  wire  T_7754;
  wire  T_7756;
  wire  T_7757;
  wire  T_7758;
  wire  T_7760;
  wire  T_7761;
  wire  T_7762;
  wire  T_7763;
  wire  fp_data_hazard_wb;
  wire  T_7764;
  wire  T_7765;
  wire  id_wb_hazard;
  reg  dcache_blocked;
  reg [31:0] GEN_408;
  wire  T_7769;
  wire  T_7770;
  reg  rocc_blocked;
  reg [31:0] GEN_409;
  wire  T_7773;
  wire  T_7776;
  wire  T_7777;
  wire  T_7778;
  wire  T_7779;
  wire  T_7780;
  wire  T_7781;
  wire  T_7784;
  wire  T_7785;
  wire  T_7786;
  wire  T_7787;
  wire  T_7788;
  wire  ctrl_stalld;
  wire  T_7790;
  wire  T_7791;
  wire  T_7792;
  wire  T_7793;
  wire  T_7794;
  wire  T_7797;
  wire [31:0] T_7798;
  wire [31:0] T_7799;
  wire  T_7800;
  wire  T_7802;
  wire  T_7803;
  wire  T_7805;
  wire  T_7806;
  wire  T_7807;
  wire  T_7810;
  wire  T_7811;
  wire  T_7812;
  wire  T_7815;
  wire  T_7816;
  wire [4:0] T_7817;
  wire [4:0] T_7820;
  wire  T_7821;
  wire  T_7822;
  wire  T_7823;
  wire  T_7826;
  wire  T_7827;
  wire  T_7830;
  wire  T_7833;
  wire  T_7834;
  wire  T_7835;
  wire  T_7838;
  wire  T_7839;
  wire  T_7840;
  wire [5:0] ex_dcache_tag;
  wire [63:0] T_7843;
  wire  T_7846;
  wire  T_7847;
  wire  T_7850;
  wire [6:0] T_7869_funct;
  wire [4:0] T_7869_rs2;
  wire [4:0] T_7869_rs1;
  wire  T_7869_xd;
  wire  T_7869_xs1;
  wire  T_7869_xs2;
  wire [4:0] T_7869_rd;
  wire [6:0] T_7869_opcode;
  wire [31:0] T_7879;
  wire [6:0] T_7880;
  wire [4:0] T_7881;
  wire  T_7882;
  wire  T_7883;
  wire  T_7884;
  wire [4:0] T_7885;
  wire [4:0] T_7886;
  wire [6:0] T_7887;
  wire [31:0] T_7888;
  wire [7:0] T_7890;
  wire [4:0] T_7891;
  reg [31:0] T_7892;
  reg [31:0] GEN_410;
  reg [31:0] T_7893;
  reg [31:0] GEN_411;
  wire [4:0] T_7894;
  reg [31:0] T_7895;
  reg [31:0] GEN_412;
  reg [31:0] T_7896;
  reg [31:0] GEN_413;
  wire  T_7898;
  reg  GEN_154;
  reg [31:0] GEN_414;
  reg [31:0] GEN_155;
  reg [31:0] GEN_415;
  reg  GEN_156;
  reg [31:0] GEN_416;
  reg [4:0] GEN_157;
  reg [31:0] GEN_417;
  reg  GEN_158;
  reg [31:0] GEN_418;
  reg  GEN_161;
  reg [31:0] GEN_419;
  reg  GEN_162;
  reg [31:0] GEN_420;
  reg  GEN_164;
  reg [31:0] GEN_421;
  reg  GEN_165;
  reg [31:0] GEN_422;
  reg  GEN_174;
  reg [31:0] GEN_423;
  reg  GEN_175;
  reg [31:0] GEN_424;
  reg  GEN_176;
  reg [31:0] GEN_425;
  reg  GEN_177;
  reg [31:0] GEN_426;
  reg  GEN_178;
  reg [31:0] GEN_427;
  reg  GEN_179;
  reg [31:0] GEN_428;
  reg  GEN_180;
  reg [31:0] GEN_429;
  reg  GEN_181;
  reg [31:0] GEN_430;
  reg  GEN_182;
  reg [31:0] GEN_431;
  reg  GEN_183;
  reg [31:0] GEN_432;
  reg  GEN_184;
  reg [31:0] GEN_433;
  reg [2:0] GEN_185;
  reg [31:0] GEN_434;
  reg [1:0] GEN_186;
  reg [31:0] GEN_435;
  reg [64:0] GEN_187;
  reg [95:0] GEN_436;
  reg [64:0] GEN_188;
  reg [95:0] GEN_437;
  reg [64:0] GEN_189;
  reg [95:0] GEN_438;
  reg  GEN_190;
  reg [31:0] GEN_439;
  reg  GEN_191;
  reg [31:0] GEN_440;
  reg  GEN_192;
  reg [31:0] GEN_441;
  reg  GEN_193;
  reg [31:0] GEN_442;
  reg  GEN_194;
  reg [31:0] GEN_443;
  reg [31:0] GEN_195;
  reg [31:0] GEN_444;
  reg [8:0] GEN_196;
  reg [31:0] GEN_445;
  reg [4:0] GEN_197;
  reg [31:0] GEN_446;
  reg [2:0] GEN_198;
  reg [31:0] GEN_447;
  reg [31:0] GEN_199;
  reg [31:0] GEN_448;
  reg  GEN_200;
  reg [31:0] GEN_449;
  reg  GEN_201;
  reg [31:0] GEN_450;
  reg [31:0] GEN_202;
  reg [31:0] GEN_451;
  reg [31:0] GEN_203;
  reg [31:0] GEN_452;
  reg  GEN_204;
  reg [31:0] GEN_453;
  reg  GEN_205;
  reg [31:0] GEN_454;
  reg  GEN_206;
  reg [31:0] GEN_455;
  reg  GEN_207;
  reg [31:0] GEN_456;
  reg  GEN_208;
  reg [31:0] GEN_457;
  reg  GEN_209;
  reg [31:0] GEN_458;
  reg  GEN_210;
  reg [31:0] GEN_459;
  reg  GEN_211;
  reg [31:0] GEN_460;
  reg [2:0] GEN_212;
  reg [31:0] GEN_461;
  reg  GEN_213;
  reg [31:0] GEN_462;
  reg [1:0] GEN_214;
  reg [31:0] GEN_463;
  reg  GEN_215;
  reg [31:0] GEN_464;
  reg [3:0] GEN_216;
  reg [31:0] GEN_465;
  reg [63:0] GEN_217;
  reg [63:0] GEN_466;
  reg  GEN_218;
  reg [31:0] GEN_467;
  reg  GEN_219;
  reg [31:0] GEN_468;
  reg [64:0] GEN_220;
  reg [95:0] GEN_469;
  reg [4:0] GEN_221;
  reg [31:0] GEN_470;
  reg  GEN_222;
  reg [31:0] GEN_471;
  reg  GEN_223;
  reg [31:0] GEN_472;
  reg  GEN_224;
  reg [31:0] GEN_473;
  reg [4:0] GEN_225;
  reg [31:0] GEN_474;
  reg [31:0] GEN_226;
  reg [31:0] GEN_475;
  reg  GEN_227;
  reg [31:0] GEN_476;
  reg [31:0] GEN_228;
  reg [31:0] GEN_477;
  reg [8:0] GEN_229;
  reg [31:0] GEN_478;
  reg [4:0] GEN_230;
  reg [31:0] GEN_479;
  reg [2:0] GEN_231;
  reg [31:0] GEN_480;
  reg  GEN_232;
  reg [31:0] GEN_481;
  reg [31:0] GEN_233;
  reg [31:0] GEN_482;
  reg  GEN_234;
  reg [31:0] GEN_483;
  reg [31:0] GEN_235;
  reg [31:0] GEN_484;
  reg  GEN_236;
  reg [31:0] GEN_485;
  reg  GEN_237;
  reg [31:0] GEN_486;
  reg  GEN_238;
  reg [31:0] GEN_487;
  reg [25:0] GEN_239;
  reg [31:0] GEN_488;
  reg  GEN_240;
  reg [31:0] GEN_489;
  reg [2:0] GEN_241;
  reg [31:0] GEN_490;
  reg  GEN_242;
  reg [31:0] GEN_491;
  reg [2:0] GEN_243;
  reg [31:0] GEN_492;
  reg [11:0] GEN_244;
  reg [31:0] GEN_493;
  reg [63:0] GEN_245;
  reg [63:0] GEN_494;
  reg  GEN_246;
  reg [31:0] GEN_495;
  reg  GEN_247;
  reg [31:0] GEN_496;
  reg [4:0] GEN_248;
  reg [31:0] GEN_497;
  reg  GEN_249;
  reg [31:0] GEN_498;
  reg  GEN_250;
  reg [31:0] GEN_499;
  reg  GEN_251;
  reg [31:0] GEN_500;
  reg  GEN_252;
  reg [31:0] GEN_501;
  reg  GEN_253;
  reg [31:0] GEN_502;
  reg  GEN_254;
  reg [31:0] GEN_503;
  reg  GEN_255;
  reg [31:0] GEN_504;
  reg  GEN_256;
  reg [31:0] GEN_505;
  reg  GEN_257;
  reg [31:0] GEN_506;
  reg  GEN_258;
  reg [31:0] GEN_507;
  reg  GEN_259;
  reg [31:0] GEN_508;
  reg  GEN_260;
  reg [31:0] GEN_509;
  reg  GEN_261;
  reg [31:0] GEN_510;
  reg  GEN_262;
  reg [31:0] GEN_511;
  reg  GEN_263;
  reg [31:0] GEN_512;
  reg  GEN_264;
  reg [31:0] GEN_513;
  reg [2:0] GEN_265;
  reg [31:0] GEN_514;
  reg [1:0] GEN_266;
  reg [31:0] GEN_515;
  reg [64:0] GEN_267;
  reg [95:0] GEN_516;
  reg [64:0] GEN_268;
  reg [95:0] GEN_517;
  reg [64:0] GEN_269;
  reg [95:0] GEN_518;
  reg  GEN_270;
  reg [31:0] GEN_519;
  CSRFile csr (
    .clk(csr_clk),
    .reset(csr_reset),
    .io_prci_reset(csr_io_prci_reset),
    .io_prci_id(csr_io_prci_id),
    .io_prci_interrupts_meip(csr_io_prci_interrupts_meip),
    .io_prci_interrupts_seip(csr_io_prci_interrupts_seip),
    .io_prci_interrupts_debug(csr_io_prci_interrupts_debug),
    .io_prci_interrupts_mtip(csr_io_prci_interrupts_mtip),
    .io_prci_interrupts_msip(csr_io_prci_interrupts_msip),
    .io_rw_addr(csr_io_rw_addr),
    .io_rw_cmd(csr_io_rw_cmd),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_wdata(csr_io_rw_wdata),
    .io_csr_stall(csr_io_csr_stall),
    .io_csr_xcpt(csr_io_csr_xcpt),
    .io_eret(csr_io_eret),
    .io_singleStep(csr_io_singleStep),
    .io_status_debug(csr_io_status_debug),
    .io_status_prv(csr_io_status_prv),
    .io_status_sd(csr_io_status_sd),
    .io_status_zero3(csr_io_status_zero3),
    .io_status_sd_rv32(csr_io_status_sd_rv32),
    .io_status_zero2(csr_io_status_zero2),
    .io_status_vm(csr_io_status_vm),
    .io_status_zero1(csr_io_status_zero1),
    .io_status_mxr(csr_io_status_mxr),
    .io_status_pum(csr_io_status_pum),
    .io_status_mprv(csr_io_status_mprv),
    .io_status_xs(csr_io_status_xs),
    .io_status_fs(csr_io_status_fs),
    .io_status_mpp(csr_io_status_mpp),
    .io_status_hpp(csr_io_status_hpp),
    .io_status_spp(csr_io_status_spp),
    .io_status_mpie(csr_io_status_mpie),
    .io_status_hpie(csr_io_status_hpie),
    .io_status_spie(csr_io_status_spie),
    .io_status_upie(csr_io_status_upie),
    .io_status_mie(csr_io_status_mie),
    .io_status_hie(csr_io_status_hie),
    .io_status_sie(csr_io_status_sie),
    .io_status_uie(csr_io_status_uie),
    .io_ptbr_asid(csr_io_ptbr_asid),
    .io_ptbr_ppn(csr_io_ptbr_ppn),
    .io_evec(csr_io_evec),
    .io_exception(csr_io_exception),
    .io_retire(csr_io_retire),
    .io_cause(csr_io_cause),
    .io_pc(csr_io_pc),
    .io_badaddr(csr_io_badaddr),
    .io_fatc(csr_io_fatc),
    .io_time(csr_io_time),
    .io_fcsr_rm(csr_io_fcsr_rm),
    .io_fcsr_flags_valid(csr_io_fcsr_flags_valid),
    .io_fcsr_flags_bits(csr_io_fcsr_flags_bits),
    .io_rocc_cmd_ready(csr_io_rocc_cmd_ready),
    .io_rocc_cmd_valid(csr_io_rocc_cmd_valid),
    .io_rocc_cmd_bits_inst_funct(csr_io_rocc_cmd_bits_inst_funct),
    .io_rocc_cmd_bits_inst_rs2(csr_io_rocc_cmd_bits_inst_rs2),
    .io_rocc_cmd_bits_inst_rs1(csr_io_rocc_cmd_bits_inst_rs1),
    .io_rocc_cmd_bits_inst_xd(csr_io_rocc_cmd_bits_inst_xd),
    .io_rocc_cmd_bits_inst_xs1(csr_io_rocc_cmd_bits_inst_xs1),
    .io_rocc_cmd_bits_inst_xs2(csr_io_rocc_cmd_bits_inst_xs2),
    .io_rocc_cmd_bits_inst_rd(csr_io_rocc_cmd_bits_inst_rd),
    .io_rocc_cmd_bits_inst_opcode(csr_io_rocc_cmd_bits_inst_opcode),
    .io_rocc_cmd_bits_rs1(csr_io_rocc_cmd_bits_rs1),
    .io_rocc_cmd_bits_rs2(csr_io_rocc_cmd_bits_rs2),
    .io_rocc_cmd_bits_status_debug(csr_io_rocc_cmd_bits_status_debug),
    .io_rocc_cmd_bits_status_prv(csr_io_rocc_cmd_bits_status_prv),
    .io_rocc_cmd_bits_status_sd(csr_io_rocc_cmd_bits_status_sd),
    .io_rocc_cmd_bits_status_zero3(csr_io_rocc_cmd_bits_status_zero3),
    .io_rocc_cmd_bits_status_sd_rv32(csr_io_rocc_cmd_bits_status_sd_rv32),
    .io_rocc_cmd_bits_status_zero2(csr_io_rocc_cmd_bits_status_zero2),
    .io_rocc_cmd_bits_status_vm(csr_io_rocc_cmd_bits_status_vm),
    .io_rocc_cmd_bits_status_zero1(csr_io_rocc_cmd_bits_status_zero1),
    .io_rocc_cmd_bits_status_mxr(csr_io_rocc_cmd_bits_status_mxr),
    .io_rocc_cmd_bits_status_pum(csr_io_rocc_cmd_bits_status_pum),
    .io_rocc_cmd_bits_status_mprv(csr_io_rocc_cmd_bits_status_mprv),
    .io_rocc_cmd_bits_status_xs(csr_io_rocc_cmd_bits_status_xs),
    .io_rocc_cmd_bits_status_fs(csr_io_rocc_cmd_bits_status_fs),
    .io_rocc_cmd_bits_status_mpp(csr_io_rocc_cmd_bits_status_mpp),
    .io_rocc_cmd_bits_status_hpp(csr_io_rocc_cmd_bits_status_hpp),
    .io_rocc_cmd_bits_status_spp(csr_io_rocc_cmd_bits_status_spp),
    .io_rocc_cmd_bits_status_mpie(csr_io_rocc_cmd_bits_status_mpie),
    .io_rocc_cmd_bits_status_hpie(csr_io_rocc_cmd_bits_status_hpie),
    .io_rocc_cmd_bits_status_spie(csr_io_rocc_cmd_bits_status_spie),
    .io_rocc_cmd_bits_status_upie(csr_io_rocc_cmd_bits_status_upie),
    .io_rocc_cmd_bits_status_mie(csr_io_rocc_cmd_bits_status_mie),
    .io_rocc_cmd_bits_status_hie(csr_io_rocc_cmd_bits_status_hie),
    .io_rocc_cmd_bits_status_sie(csr_io_rocc_cmd_bits_status_sie),
    .io_rocc_cmd_bits_status_uie(csr_io_rocc_cmd_bits_status_uie),
    .io_rocc_resp_ready(csr_io_rocc_resp_ready),
    .io_rocc_resp_valid(csr_io_rocc_resp_valid),
    .io_rocc_resp_bits_rd(csr_io_rocc_resp_bits_rd),
    .io_rocc_resp_bits_data(csr_io_rocc_resp_bits_data),
    .io_rocc_mem_req_ready(csr_io_rocc_mem_req_ready),
    .io_rocc_mem_req_valid(csr_io_rocc_mem_req_valid),
    .io_rocc_mem_req_bits_addr(csr_io_rocc_mem_req_bits_addr),
    .io_rocc_mem_req_bits_tag(csr_io_rocc_mem_req_bits_tag),
    .io_rocc_mem_req_bits_cmd(csr_io_rocc_mem_req_bits_cmd),
    .io_rocc_mem_req_bits_typ(csr_io_rocc_mem_req_bits_typ),
    .io_rocc_mem_req_bits_phys(csr_io_rocc_mem_req_bits_phys),
    .io_rocc_mem_req_bits_data(csr_io_rocc_mem_req_bits_data),
    .io_rocc_mem_s1_kill(csr_io_rocc_mem_s1_kill),
    .io_rocc_mem_s1_data(csr_io_rocc_mem_s1_data),
    .io_rocc_mem_s2_nack(csr_io_rocc_mem_s2_nack),
    .io_rocc_mem_resp_valid(csr_io_rocc_mem_resp_valid),
    .io_rocc_mem_resp_bits_addr(csr_io_rocc_mem_resp_bits_addr),
    .io_rocc_mem_resp_bits_tag(csr_io_rocc_mem_resp_bits_tag),
    .io_rocc_mem_resp_bits_cmd(csr_io_rocc_mem_resp_bits_cmd),
    .io_rocc_mem_resp_bits_typ(csr_io_rocc_mem_resp_bits_typ),
    .io_rocc_mem_resp_bits_data(csr_io_rocc_mem_resp_bits_data),
    .io_rocc_mem_resp_bits_replay(csr_io_rocc_mem_resp_bits_replay),
    .io_rocc_mem_resp_bits_has_data(csr_io_rocc_mem_resp_bits_has_data),
    .io_rocc_mem_resp_bits_data_word_bypass(csr_io_rocc_mem_resp_bits_data_word_bypass),
    .io_rocc_mem_resp_bits_store_data(csr_io_rocc_mem_resp_bits_store_data),
    .io_rocc_mem_replay_next(csr_io_rocc_mem_replay_next),
    .io_rocc_mem_xcpt_ma_ld(csr_io_rocc_mem_xcpt_ma_ld),
    .io_rocc_mem_xcpt_ma_st(csr_io_rocc_mem_xcpt_ma_st),
    .io_rocc_mem_xcpt_pf_ld(csr_io_rocc_mem_xcpt_pf_ld),
    .io_rocc_mem_xcpt_pf_st(csr_io_rocc_mem_xcpt_pf_st),
    .io_rocc_mem_invalidate_lr(csr_io_rocc_mem_invalidate_lr),
    .io_rocc_mem_ordered(csr_io_rocc_mem_ordered),
    .io_rocc_busy(csr_io_rocc_busy),
    .io_rocc_interrupt(csr_io_rocc_interrupt),
    .io_rocc_autl_acquire_ready(csr_io_rocc_autl_acquire_ready),
    .io_rocc_autl_acquire_valid(csr_io_rocc_autl_acquire_valid),
    .io_rocc_autl_acquire_bits_addr_block(csr_io_rocc_autl_acquire_bits_addr_block),
    .io_rocc_autl_acquire_bits_client_xact_id(csr_io_rocc_autl_acquire_bits_client_xact_id),
    .io_rocc_autl_acquire_bits_addr_beat(csr_io_rocc_autl_acquire_bits_addr_beat),
    .io_rocc_autl_acquire_bits_is_builtin_type(csr_io_rocc_autl_acquire_bits_is_builtin_type),
    .io_rocc_autl_acquire_bits_a_type(csr_io_rocc_autl_acquire_bits_a_type),
    .io_rocc_autl_acquire_bits_union(csr_io_rocc_autl_acquire_bits_union),
    .io_rocc_autl_acquire_bits_data(csr_io_rocc_autl_acquire_bits_data),
    .io_rocc_autl_grant_ready(csr_io_rocc_autl_grant_ready),
    .io_rocc_autl_grant_valid(csr_io_rocc_autl_grant_valid),
    .io_rocc_autl_grant_bits_addr_beat(csr_io_rocc_autl_grant_bits_addr_beat),
    .io_rocc_autl_grant_bits_client_xact_id(csr_io_rocc_autl_grant_bits_client_xact_id),
    .io_rocc_autl_grant_bits_manager_xact_id(csr_io_rocc_autl_grant_bits_manager_xact_id),
    .io_rocc_autl_grant_bits_is_builtin_type(csr_io_rocc_autl_grant_bits_is_builtin_type),
    .io_rocc_autl_grant_bits_g_type(csr_io_rocc_autl_grant_bits_g_type),
    .io_rocc_autl_grant_bits_data(csr_io_rocc_autl_grant_bits_data),
    .io_rocc_fpu_req_ready(csr_io_rocc_fpu_req_ready),
    .io_rocc_fpu_req_valid(csr_io_rocc_fpu_req_valid),
    .io_rocc_fpu_req_bits_cmd(csr_io_rocc_fpu_req_bits_cmd),
    .io_rocc_fpu_req_bits_ldst(csr_io_rocc_fpu_req_bits_ldst),
    .io_rocc_fpu_req_bits_wen(csr_io_rocc_fpu_req_bits_wen),
    .io_rocc_fpu_req_bits_ren1(csr_io_rocc_fpu_req_bits_ren1),
    .io_rocc_fpu_req_bits_ren2(csr_io_rocc_fpu_req_bits_ren2),
    .io_rocc_fpu_req_bits_ren3(csr_io_rocc_fpu_req_bits_ren3),
    .io_rocc_fpu_req_bits_swap12(csr_io_rocc_fpu_req_bits_swap12),
    .io_rocc_fpu_req_bits_swap23(csr_io_rocc_fpu_req_bits_swap23),
    .io_rocc_fpu_req_bits_single(csr_io_rocc_fpu_req_bits_single),
    .io_rocc_fpu_req_bits_fromint(csr_io_rocc_fpu_req_bits_fromint),
    .io_rocc_fpu_req_bits_toint(csr_io_rocc_fpu_req_bits_toint),
    .io_rocc_fpu_req_bits_fastpipe(csr_io_rocc_fpu_req_bits_fastpipe),
    .io_rocc_fpu_req_bits_fma(csr_io_rocc_fpu_req_bits_fma),
    .io_rocc_fpu_req_bits_div(csr_io_rocc_fpu_req_bits_div),
    .io_rocc_fpu_req_bits_sqrt(csr_io_rocc_fpu_req_bits_sqrt),
    .io_rocc_fpu_req_bits_round(csr_io_rocc_fpu_req_bits_round),
    .io_rocc_fpu_req_bits_wflags(csr_io_rocc_fpu_req_bits_wflags),
    .io_rocc_fpu_req_bits_rm(csr_io_rocc_fpu_req_bits_rm),
    .io_rocc_fpu_req_bits_typ(csr_io_rocc_fpu_req_bits_typ),
    .io_rocc_fpu_req_bits_in1(csr_io_rocc_fpu_req_bits_in1),
    .io_rocc_fpu_req_bits_in2(csr_io_rocc_fpu_req_bits_in2),
    .io_rocc_fpu_req_bits_in3(csr_io_rocc_fpu_req_bits_in3),
    .io_rocc_fpu_resp_ready(csr_io_rocc_fpu_resp_ready),
    .io_rocc_fpu_resp_valid(csr_io_rocc_fpu_resp_valid),
    .io_rocc_fpu_resp_bits_data(csr_io_rocc_fpu_resp_bits_data),
    .io_rocc_fpu_resp_bits_exc(csr_io_rocc_fpu_resp_bits_exc),
    .io_rocc_exception(csr_io_rocc_exception),
    .io_rocc_csr_waddr(csr_io_rocc_csr_waddr),
    .io_rocc_csr_wdata(csr_io_rocc_csr_wdata),
    .io_rocc_csr_wen(csr_io_rocc_csr_wen),
    .io_rocc_host_id(csr_io_rocc_host_id),
    .io_interrupt(csr_io_interrupt),
    .io_interrupt_cause(csr_io_interrupt_cause),
    .io_bp_0_control_tdrtype(csr_io_bp_0_control_tdrtype),
    .io_bp_0_control_bpamaskmax(csr_io_bp_0_control_bpamaskmax),
    .io_bp_0_control_reserved(csr_io_bp_0_control_reserved),
    .io_bp_0_control_bpaction(csr_io_bp_0_control_bpaction),
    .io_bp_0_control_bpmatch(csr_io_bp_0_control_bpmatch),
    .io_bp_0_control_m(csr_io_bp_0_control_m),
    .io_bp_0_control_h(csr_io_bp_0_control_h),
    .io_bp_0_control_s(csr_io_bp_0_control_s),
    .io_bp_0_control_u(csr_io_bp_0_control_u),
    .io_bp_0_control_r(csr_io_bp_0_control_r),
    .io_bp_0_control_w(csr_io_bp_0_control_w),
    .io_bp_0_control_x(csr_io_bp_0_control_x),
    .io_bp_0_address(csr_io_bp_0_address),
    .io_bp_1_control_tdrtype(csr_io_bp_1_control_tdrtype),
    .io_bp_1_control_bpamaskmax(csr_io_bp_1_control_bpamaskmax),
    .io_bp_1_control_reserved(csr_io_bp_1_control_reserved),
    .io_bp_1_control_bpaction(csr_io_bp_1_control_bpaction),
    .io_bp_1_control_bpmatch(csr_io_bp_1_control_bpmatch),
    .io_bp_1_control_m(csr_io_bp_1_control_m),
    .io_bp_1_control_h(csr_io_bp_1_control_h),
    .io_bp_1_control_s(csr_io_bp_1_control_s),
    .io_bp_1_control_u(csr_io_bp_1_control_u),
    .io_bp_1_control_r(csr_io_bp_1_control_r),
    .io_bp_1_control_w(csr_io_bp_1_control_w),
    .io_bp_1_control_x(csr_io_bp_1_control_x),
    .io_bp_1_address(csr_io_bp_1_address)
  );
  BreakpointUnit bpu (
    .clk(bpu_clk),
    .reset(bpu_reset),
    .io_status_debug(bpu_io_status_debug),
    .io_status_prv(bpu_io_status_prv),
    .io_status_sd(bpu_io_status_sd),
    .io_status_zero3(bpu_io_status_zero3),
    .io_status_sd_rv32(bpu_io_status_sd_rv32),
    .io_status_zero2(bpu_io_status_zero2),
    .io_status_vm(bpu_io_status_vm),
    .io_status_zero1(bpu_io_status_zero1),
    .io_status_mxr(bpu_io_status_mxr),
    .io_status_pum(bpu_io_status_pum),
    .io_status_mprv(bpu_io_status_mprv),
    .io_status_xs(bpu_io_status_xs),
    .io_status_fs(bpu_io_status_fs),
    .io_status_mpp(bpu_io_status_mpp),
    .io_status_hpp(bpu_io_status_hpp),
    .io_status_spp(bpu_io_status_spp),
    .io_status_mpie(bpu_io_status_mpie),
    .io_status_hpie(bpu_io_status_hpie),
    .io_status_spie(bpu_io_status_spie),
    .io_status_upie(bpu_io_status_upie),
    .io_status_mie(bpu_io_status_mie),
    .io_status_hie(bpu_io_status_hie),
    .io_status_sie(bpu_io_status_sie),
    .io_status_uie(bpu_io_status_uie),
    .io_bp_0_control_tdrtype(bpu_io_bp_0_control_tdrtype),
    .io_bp_0_control_bpamaskmax(bpu_io_bp_0_control_bpamaskmax),
    .io_bp_0_control_reserved(bpu_io_bp_0_control_reserved),
    .io_bp_0_control_bpaction(bpu_io_bp_0_control_bpaction),
    .io_bp_0_control_bpmatch(bpu_io_bp_0_control_bpmatch),
    .io_bp_0_control_m(bpu_io_bp_0_control_m),
    .io_bp_0_control_h(bpu_io_bp_0_control_h),
    .io_bp_0_control_s(bpu_io_bp_0_control_s),
    .io_bp_0_control_u(bpu_io_bp_0_control_u),
    .io_bp_0_control_r(bpu_io_bp_0_control_r),
    .io_bp_0_control_w(bpu_io_bp_0_control_w),
    .io_bp_0_control_x(bpu_io_bp_0_control_x),
    .io_bp_0_address(bpu_io_bp_0_address),
    .io_bp_1_control_tdrtype(bpu_io_bp_1_control_tdrtype),
    .io_bp_1_control_bpamaskmax(bpu_io_bp_1_control_bpamaskmax),
    .io_bp_1_control_reserved(bpu_io_bp_1_control_reserved),
    .io_bp_1_control_bpaction(bpu_io_bp_1_control_bpaction),
    .io_bp_1_control_bpmatch(bpu_io_bp_1_control_bpmatch),
    .io_bp_1_control_m(bpu_io_bp_1_control_m),
    .io_bp_1_control_h(bpu_io_bp_1_control_h),
    .io_bp_1_control_s(bpu_io_bp_1_control_s),
    .io_bp_1_control_u(bpu_io_bp_1_control_u),
    .io_bp_1_control_r(bpu_io_bp_1_control_r),
    .io_bp_1_control_w(bpu_io_bp_1_control_w),
    .io_bp_1_control_x(bpu_io_bp_1_control_x),
    .io_bp_1_address(bpu_io_bp_1_address),
    .io_pc(bpu_io_pc),
    .io_ea(bpu_io_ea),
    .io_xcpt_if(bpu_io_xcpt_if),
    .io_xcpt_ld(bpu_io_xcpt_ld),
    .io_xcpt_st(bpu_io_xcpt_st)
  );
  ALU alu (
    .clk(alu_clk),
    .reset(alu_reset),
    .io_dw(alu_io_dw),
    .io_fn(alu_io_fn),
    .io_in2(alu_io_in2),
    .io_in1(alu_io_in1),
    .io_out(alu_io_out),
    .io_adder_out(alu_io_adder_out),
    .io_cmp_out(alu_io_cmp_out)
  );
  MulDiv div (
    .clk(div_clk),
    .reset(div_reset),
    .io_req_ready(div_io_req_ready),
    .io_req_valid(div_io_req_valid),
    .io_req_bits_fn(div_io_req_bits_fn),
    .io_req_bits_dw(div_io_req_bits_dw),
    .io_req_bits_in1(div_io_req_bits_in1),
    .io_req_bits_in2(div_io_req_bits_in2),
    .io_req_bits_tag(div_io_req_bits_tag),
    .io_kill(div_io_kill),
    .io_resp_ready(div_io_resp_ready),
    .io_resp_valid(div_io_resp_valid),
    .io_resp_bits_data(div_io_resp_bits_data),
    .io_resp_bits_tag(div_io_resp_bits_tag)
  );
  assign io_imem_req_valid = take_pc_mem_wb;
  assign io_imem_req_bits_pc = T_7799;
  assign io_imem_req_bits_speculative = T_7604;
  assign io_imem_resp_ready = T_7807;
  assign io_imem_btb_update_valid = T_7815;
  assign io_imem_btb_update_bits_prediction_valid = mem_reg_btb_hit;
  assign io_imem_btb_update_bits_prediction_bits_taken = mem_reg_btb_resp_taken;
  assign io_imem_btb_update_bits_prediction_bits_mask = mem_reg_btb_resp_mask;
  assign io_imem_btb_update_bits_prediction_bits_bridx = mem_reg_btb_resp_bridx;
  assign io_imem_btb_update_bits_prediction_bits_target = mem_reg_btb_resp_target;
  assign io_imem_btb_update_bits_prediction_bits_entry = mem_reg_btb_resp_entry;
  assign io_imem_btb_update_bits_prediction_bits_bht_history = mem_reg_btb_resp_bht_history;
  assign io_imem_btb_update_bits_prediction_bits_bht_value = mem_reg_btb_resp_bht_value;
  assign io_imem_btb_update_bits_pc = mem_reg_pc;
  assign io_imem_btb_update_bits_target = io_imem_req_bits_pc;
  assign io_imem_btb_update_bits_taken = GEN_154;
  assign io_imem_btb_update_bits_isJump = T_7816;
  assign io_imem_btb_update_bits_isReturn = T_7822;
  assign io_imem_btb_update_bits_br_pc = mem_reg_pc;
  assign io_imem_bht_update_valid = T_7826;
  assign io_imem_bht_update_bits_prediction_valid = io_imem_btb_update_bits_prediction_valid;
  assign io_imem_bht_update_bits_prediction_bits_taken = io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_bht_update_bits_prediction_bits_mask = io_imem_btb_update_bits_prediction_bits_mask;
  assign io_imem_bht_update_bits_prediction_bits_bridx = io_imem_btb_update_bits_prediction_bits_bridx;
  assign io_imem_bht_update_bits_prediction_bits_target = io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_bht_update_bits_prediction_bits_entry = io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_bht_update_bits_prediction_bits_bht_history = io_imem_btb_update_bits_prediction_bits_bht_history;
  assign io_imem_bht_update_bits_prediction_bits_bht_value = io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_bht_update_bits_pc = mem_reg_pc;
  assign io_imem_bht_update_bits_taken = mem_br_taken;
  assign io_imem_bht_update_bits_mispredict = mem_wrong_npc;
  assign io_imem_ras_update_valid = T_7833;
  assign io_imem_ras_update_bits_isCall = T_7835;
  assign io_imem_ras_update_bits_isReturn = io_imem_btb_update_bits_isReturn;
  assign io_imem_ras_update_bits_returnAddr = mem_int_wdata;
  assign io_imem_ras_update_bits_prediction_valid = io_imem_btb_update_bits_prediction_valid;
  assign io_imem_ras_update_bits_prediction_bits_taken = io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_ras_update_bits_prediction_bits_mask = io_imem_btb_update_bits_prediction_bits_mask;
  assign io_imem_ras_update_bits_prediction_bits_bridx = io_imem_btb_update_bits_prediction_bits_bridx;
  assign io_imem_ras_update_bits_prediction_bits_target = io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_ras_update_bits_prediction_bits_entry = io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_ras_update_bits_prediction_bits_bht_history = io_imem_btb_update_bits_prediction_bits_bht_history;
  assign io_imem_ras_update_bits_prediction_bits_bht_value = io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_flush_icache = T_7803;
  assign io_imem_flush_tlb = csr_io_fatc;
  assign io_dmem_req_valid = T_7840;
  assign io_dmem_req_bits_addr = alu_io_adder_out;
  assign io_dmem_req_bits_tag = {{3'd0}, ex_dcache_tag};
  assign io_dmem_req_bits_cmd = ex_ctrl_mem_cmd;
  assign io_dmem_req_bits_typ = ex_ctrl_mem_type;
  assign io_dmem_req_bits_phys = 1'h0;
  assign io_dmem_req_bits_data = GEN_155;
  assign io_dmem_s1_kill = T_7600;
  assign io_dmem_s1_data = T_7843[31:0];
  assign io_dmem_invalidate_lr = wb_xcpt;
  assign io_ptw_ptbr_asid = csr_io_ptbr_asid;
  assign io_ptw_ptbr_ppn = csr_io_ptbr_ppn;
  assign io_ptw_invalidate = csr_io_fatc;
  assign io_ptw_status_debug = csr_io_status_debug;
  assign io_ptw_status_prv = csr_io_status_prv;
  assign io_ptw_status_sd = csr_io_status_sd;
  assign io_ptw_status_zero3 = csr_io_status_zero3;
  assign io_ptw_status_sd_rv32 = csr_io_status_sd_rv32;
  assign io_ptw_status_zero2 = csr_io_status_zero2;
  assign io_ptw_status_vm = csr_io_status_vm;
  assign io_ptw_status_zero1 = csr_io_status_zero1;
  assign io_ptw_status_mxr = csr_io_status_mxr;
  assign io_ptw_status_pum = csr_io_status_pum;
  assign io_ptw_status_mprv = csr_io_status_mprv;
  assign io_ptw_status_xs = csr_io_status_xs;
  assign io_ptw_status_fs = csr_io_status_fs;
  assign io_ptw_status_mpp = csr_io_status_mpp;
  assign io_ptw_status_hpp = csr_io_status_hpp;
  assign io_ptw_status_spp = csr_io_status_spp;
  assign io_ptw_status_mpie = csr_io_status_mpie;
  assign io_ptw_status_hpie = csr_io_status_hpie;
  assign io_ptw_status_spie = csr_io_status_spie;
  assign io_ptw_status_upie = csr_io_status_upie;
  assign io_ptw_status_mie = csr_io_status_mie;
  assign io_ptw_status_hie = csr_io_status_hie;
  assign io_ptw_status_sie = csr_io_status_sie;
  assign io_ptw_status_uie = csr_io_status_uie;
  assign io_fpu_inst = io_imem_resp_bits_data_0;
  assign io_fpu_fromint_data = T_7191;
  assign io_fpu_fcsr_rm = csr_io_fcsr_rm;
  assign io_fpu_dmem_resp_val = T_7839;
  assign io_fpu_dmem_resp_type = io_dmem_resp_bits_typ;
  assign io_fpu_dmem_resp_tag = dmem_resp_waddr[4:0];
  assign io_fpu_dmem_resp_data = {{32'd0}, io_dmem_resp_bits_data_word_bypass};
  assign io_fpu_valid = T_7838;
  assign io_fpu_killx = ctrl_killx;
  assign io_fpu_killm = killm_common;
  assign io_fpu_cp_req_valid = GEN_156;
  assign io_fpu_cp_req_bits_cmd = GEN_157;
  assign io_fpu_cp_req_bits_ldst = GEN_158;
  assign io_fpu_cp_req_bits_wen = GEN_161;
  assign io_fpu_cp_req_bits_ren1 = GEN_162;
  assign io_fpu_cp_req_bits_ren2 = GEN_164;
  assign io_fpu_cp_req_bits_ren3 = GEN_165;
  assign io_fpu_cp_req_bits_swap12 = GEN_174;
  assign io_fpu_cp_req_bits_swap23 = GEN_175;
  assign io_fpu_cp_req_bits_single = GEN_176;
  assign io_fpu_cp_req_bits_fromint = GEN_177;
  assign io_fpu_cp_req_bits_toint = GEN_178;
  assign io_fpu_cp_req_bits_fastpipe = GEN_179;
  assign io_fpu_cp_req_bits_fma = GEN_180;
  assign io_fpu_cp_req_bits_div = GEN_181;
  assign io_fpu_cp_req_bits_sqrt = GEN_182;
  assign io_fpu_cp_req_bits_round = GEN_183;
  assign io_fpu_cp_req_bits_wflags = GEN_184;
  assign io_fpu_cp_req_bits_rm = GEN_185;
  assign io_fpu_cp_req_bits_typ = GEN_186;
  assign io_fpu_cp_req_bits_in1 = GEN_187;
  assign io_fpu_cp_req_bits_in2 = GEN_188;
  assign io_fpu_cp_req_bits_in3 = GEN_189;
  assign io_fpu_cp_resp_ready = GEN_190;
  assign io_rocc_cmd_valid = T_7847;
  assign io_rocc_cmd_bits_inst_funct = T_7869_funct;
  assign io_rocc_cmd_bits_inst_rs2 = T_7869_rs2;
  assign io_rocc_cmd_bits_inst_rs1 = T_7869_rs1;
  assign io_rocc_cmd_bits_inst_xd = T_7869_xd;
  assign io_rocc_cmd_bits_inst_xs1 = T_7869_xs1;
  assign io_rocc_cmd_bits_inst_xs2 = T_7869_xs2;
  assign io_rocc_cmd_bits_inst_rd = T_7869_rd;
  assign io_rocc_cmd_bits_inst_opcode = T_7869_opcode;
  assign io_rocc_cmd_bits_rs1 = wb_reg_wdata;
  assign io_rocc_cmd_bits_rs2 = wb_reg_rs2;
  assign io_rocc_cmd_bits_status_debug = csr_io_status_debug;
  assign io_rocc_cmd_bits_status_prv = csr_io_status_prv;
  assign io_rocc_cmd_bits_status_sd = csr_io_status_sd;
  assign io_rocc_cmd_bits_status_zero3 = csr_io_status_zero3;
  assign io_rocc_cmd_bits_status_sd_rv32 = csr_io_status_sd_rv32;
  assign io_rocc_cmd_bits_status_zero2 = csr_io_status_zero2;
  assign io_rocc_cmd_bits_status_vm = csr_io_status_vm;
  assign io_rocc_cmd_bits_status_zero1 = csr_io_status_zero1;
  assign io_rocc_cmd_bits_status_mxr = csr_io_status_mxr;
  assign io_rocc_cmd_bits_status_pum = csr_io_status_pum;
  assign io_rocc_cmd_bits_status_mprv = csr_io_status_mprv;
  assign io_rocc_cmd_bits_status_xs = csr_io_status_xs;
  assign io_rocc_cmd_bits_status_fs = csr_io_status_fs;
  assign io_rocc_cmd_bits_status_mpp = csr_io_status_mpp;
  assign io_rocc_cmd_bits_status_hpp = csr_io_status_hpp;
  assign io_rocc_cmd_bits_status_spp = csr_io_status_spp;
  assign io_rocc_cmd_bits_status_mpie = csr_io_status_mpie;
  assign io_rocc_cmd_bits_status_hpie = csr_io_status_hpie;
  assign io_rocc_cmd_bits_status_spie = csr_io_status_spie;
  assign io_rocc_cmd_bits_status_upie = csr_io_status_upie;
  assign io_rocc_cmd_bits_status_mie = csr_io_status_mie;
  assign io_rocc_cmd_bits_status_hie = csr_io_status_hie;
  assign io_rocc_cmd_bits_status_sie = csr_io_status_sie;
  assign io_rocc_cmd_bits_status_uie = csr_io_status_uie;
  assign io_rocc_resp_ready = GEN_191;
  assign io_rocc_mem_req_ready = GEN_192;
  assign io_rocc_mem_s2_nack = GEN_193;
  assign io_rocc_mem_resp_valid = GEN_194;
  assign io_rocc_mem_resp_bits_addr = GEN_195;
  assign io_rocc_mem_resp_bits_tag = GEN_196;
  assign io_rocc_mem_resp_bits_cmd = GEN_197;
  assign io_rocc_mem_resp_bits_typ = GEN_198;
  assign io_rocc_mem_resp_bits_data = GEN_199;
  assign io_rocc_mem_resp_bits_replay = GEN_200;
  assign io_rocc_mem_resp_bits_has_data = GEN_201;
  assign io_rocc_mem_resp_bits_data_word_bypass = GEN_202;
  assign io_rocc_mem_resp_bits_store_data = GEN_203;
  assign io_rocc_mem_replay_next = GEN_204;
  assign io_rocc_mem_xcpt_ma_ld = GEN_205;
  assign io_rocc_mem_xcpt_ma_st = GEN_206;
  assign io_rocc_mem_xcpt_pf_ld = GEN_207;
  assign io_rocc_mem_xcpt_pf_st = GEN_208;
  assign io_rocc_mem_ordered = GEN_209;
  assign io_rocc_autl_acquire_ready = GEN_210;
  assign io_rocc_autl_grant_valid = GEN_211;
  assign io_rocc_autl_grant_bits_addr_beat = GEN_212;
  assign io_rocc_autl_grant_bits_client_xact_id = GEN_213;
  assign io_rocc_autl_grant_bits_manager_xact_id = GEN_214;
  assign io_rocc_autl_grant_bits_is_builtin_type = GEN_215;
  assign io_rocc_autl_grant_bits_g_type = GEN_216;
  assign io_rocc_autl_grant_bits_data = GEN_217;
  assign io_rocc_fpu_req_ready = GEN_218;
  assign io_rocc_fpu_resp_valid = GEN_219;
  assign io_rocc_fpu_resp_bits_data = GEN_220;
  assign io_rocc_fpu_resp_bits_exc = GEN_221;
  assign io_rocc_exception = T_7850;
  assign io_rocc_csr_waddr = csr_io_rocc_csr_waddr;
  assign io_rocc_csr_wdata = csr_io_rocc_csr_wdata;
  assign io_rocc_csr_wen = csr_io_rocc_csr_wen;
  assign io_rocc_host_id = GEN_222;
  assign take_pc_mem = T_7532;
  assign take_pc_wb = T_7623;
  assign take_pc_mem_wb = take_pc_wb | take_pc_mem;
  assign id_ctrl_legal = T_6660;
  assign id_ctrl_fp = 1'h0;
  assign id_ctrl_rocc = 1'h0;
  assign id_ctrl_branch = T_6666;
  assign id_ctrl_jal = T_6672;
  assign id_ctrl_jalr = T_6678;
  assign id_ctrl_rxs2 = T_6691;
  assign id_ctrl_rxs1 = T_6707;
  assign id_ctrl_sel_alu2 = T_6741;
  assign id_ctrl_sel_alu1 = T_6757;
  assign id_ctrl_sel_imm = T_6785;
  assign id_ctrl_alu_dw = 1'h1;
  assign id_ctrl_alu_fn = T_6875;
  assign id_ctrl_mem = T_6888;
  assign id_ctrl_mem_cmd = T_6904;
  assign id_ctrl_mem_type = T_6924;
  assign id_ctrl_rfs1 = 1'h0;
  assign id_ctrl_rfs2 = 1'h0;
  assign id_ctrl_rfs3 = 1'h0;
  assign id_ctrl_wfd = 1'h0;
  assign id_ctrl_div = T_6932;
  assign id_ctrl_wxd = T_6961;
  assign id_ctrl_csr = T_6981;
  assign id_ctrl_fence_i = T_6985;
  assign id_ctrl_fence = T_6991;
  assign id_ctrl_amo = 1'h0;
  assign T_6562 = io_imem_resp_bits_data_0 & 32'h505f;
  assign T_6564 = T_6562 == 32'h3;
  assign T_6566 = io_imem_resp_bits_data_0 & 32'h207f;
  assign T_6568 = T_6566 == 32'h3;
  assign T_6570 = io_imem_resp_bits_data_0 & 32'h607f;
  assign T_6572 = T_6570 == 32'hf;
  assign T_6574 = io_imem_resp_bits_data_0 & 32'h5f;
  assign T_6576 = T_6574 == 32'h17;
  assign T_6578 = io_imem_resp_bits_data_0 & 32'hfc00007f;
  assign T_6580 = T_6578 == 32'h33;
  assign T_6582 = io_imem_resp_bits_data_0 & 32'hbe00707f;
  assign T_6584 = T_6582 == 32'h33;
  assign T_6586 = io_imem_resp_bits_data_0 & 32'h707b;
  assign T_6588 = T_6586 == 32'h63;
  assign T_6590 = io_imem_resp_bits_data_0 & 32'h7f;
  assign T_6592 = T_6590 == 32'h6f;
  assign T_6594 = io_imem_resp_bits_data_0 & 32'hffefffff;
  assign T_6596 = T_6594 == 32'h73;
  assign T_6598 = io_imem_resp_bits_data_0 & 32'hfc00305f;
  assign T_6600 = T_6598 == 32'h1013;
  assign T_6604 = T_6566 == 32'h2013;
  assign T_6608 = T_6566 == 32'h2073;
  assign T_6610 = io_imem_resp_bits_data_0 & 32'hbc00707f;
  assign T_6612 = T_6610 == 32'h5013;
  assign T_6616 = T_6582 == 32'h5033;
  assign T_6618 = io_imem_resp_bits_data_0 == 32'h10500073;
  assign T_6620 = io_imem_resp_bits_data_0 == 32'h30200073;
  assign T_6622 = io_imem_resp_bits_data_0 == 32'h7b200073;
  assign T_6624 = io_imem_resp_bits_data_0 & 32'h603f;
  assign T_6626 = T_6624 == 32'h23;
  assign T_6628 = io_imem_resp_bits_data_0 & 32'h306f;
  assign T_6630 = T_6628 == 32'h1063;
  assign T_6632 = io_imem_resp_bits_data_0 & 32'h407f;
  assign T_6634 = T_6632 == 32'h4063;
  assign T_6638 = T_6628 == 32'h3;
  assign T_6641 = T_6564 | T_6568;
  assign T_6642 = T_6641 | T_6572;
  assign T_6643 = T_6642 | T_6576;
  assign T_6644 = T_6643 | T_6580;
  assign T_6645 = T_6644 | T_6584;
  assign T_6646 = T_6645 | T_6588;
  assign T_6647 = T_6646 | T_6592;
  assign T_6648 = T_6647 | T_6596;
  assign T_6649 = T_6648 | T_6600;
  assign T_6650 = T_6649 | T_6604;
  assign T_6651 = T_6650 | T_6608;
  assign T_6652 = T_6651 | T_6612;
  assign T_6653 = T_6652 | T_6616;
  assign T_6654 = T_6653 | T_6618;
  assign T_6655 = T_6654 | T_6620;
  assign T_6656 = T_6655 | T_6622;
  assign T_6657 = T_6656 | T_6626;
  assign T_6658 = T_6657 | T_6630;
  assign T_6659 = T_6658 | T_6634;
  assign T_6660 = T_6659 | T_6638;
  assign T_6664 = io_imem_resp_bits_data_0 & 32'h54;
  assign T_6666 = T_6664 == 32'h40;
  assign T_6670 = io_imem_resp_bits_data_0 & 32'h48;
  assign T_6672 = T_6670 == 32'h48;
  assign T_6676 = io_imem_resp_bits_data_0 & 32'h1c;
  assign T_6678 = T_6676 == 32'h4;
  assign T_6682 = io_imem_resp_bits_data_0 & 32'h64;
  assign T_6684 = T_6682 == 32'h20;
  assign T_6686 = io_imem_resp_bits_data_0 & 32'h34;
  assign T_6688 = T_6686 == 32'h20;
  assign T_6691 = T_6684 | T_6688;
  assign T_6693 = io_imem_resp_bits_data_0 & 32'h4004;
  assign T_6695 = T_6693 == 32'h0;
  assign T_6697 = io_imem_resp_bits_data_0 & 32'h44;
  assign T_6699 = T_6697 == 32'h0;
  assign T_6701 = io_imem_resp_bits_data_0 & 32'h18;
  assign T_6703 = T_6701 == 32'h0;
  assign T_6706 = T_6695 | T_6699;
  assign T_6707 = T_6706 | T_6703;
  assign T_6709 = io_imem_resp_bits_data_0 & 32'h50;
  assign T_6711 = T_6709 == 32'h0;
  assign T_6713 = io_imem_resp_bits_data_0 & 32'h20;
  assign T_6715 = T_6713 == 32'h0;
  assign T_6717 = io_imem_resp_bits_data_0 & 32'h4;
  assign T_6719 = T_6717 == 32'h4;
  assign T_6721 = io_imem_resp_bits_data_0 & 32'h4050;
  assign T_6723 = T_6721 == 32'h4050;
  assign T_6726 = T_6711 | T_6715;
  assign T_6727 = T_6726 | T_6719;
  assign T_6728 = T_6727 | T_6723;
  assign T_6730 = io_imem_resp_bits_data_0 & 32'h40;
  assign T_6732 = T_6730 == 32'h0;
  assign T_6734 = io_imem_resp_bits_data_0 & 32'h4008;
  assign T_6736 = T_6734 == 32'h4000;
  assign T_6739 = T_6732 | T_6703;
  assign T_6740 = T_6739 | T_6736;
  assign T_6741 = {T_6740,T_6728};
  assign T_6747 = io_imem_resp_bits_data_0 & 32'h24;
  assign T_6749 = T_6747 == 32'h4;
  assign T_6751 = io_imem_resp_bits_data_0 & 32'h8;
  assign T_6753 = T_6751 == 32'h8;
  assign T_6756 = T_6749 | T_6753;
  assign T_6757 = {T_6756,T_6707};
  assign T_6761 = T_6697 == 32'h40;
  assign T_6764 = T_6753 | T_6761;
  assign T_6768 = T_6697 == 32'h4;
  assign T_6771 = T_6768 | T_6753;
  assign T_6775 = T_6747 == 32'h0;
  assign T_6777 = io_imem_resp_bits_data_0 & 32'h14;
  assign T_6779 = T_6777 == 32'h10;
  assign T_6782 = T_6775 | T_6678;
  assign T_6783 = T_6782 | T_6779;
  assign T_6784 = {T_6771,T_6764};
  assign T_6785 = {T_6783,T_6784};
  assign T_6793 = io_imem_resp_bits_data_0 & 32'h3054;
  assign T_6795 = T_6793 == 32'h1010;
  assign T_6797 = io_imem_resp_bits_data_0 & 32'h1058;
  assign T_6799 = T_6797 == 32'h1040;
  assign T_6801 = io_imem_resp_bits_data_0 & 32'h7044;
  assign T_6803 = T_6801 == 32'h7000;
  assign T_6806 = T_6795 | T_6799;
  assign T_6807 = T_6806 | T_6803;
  assign T_6809 = io_imem_resp_bits_data_0 & 32'h4054;
  assign T_6811 = T_6809 == 32'h40;
  assign T_6813 = io_imem_resp_bits_data_0 & 32'h3044;
  assign T_6815 = T_6813 == 32'h3000;
  assign T_6817 = io_imem_resp_bits_data_0 & 32'h6044;
  assign T_6819 = T_6817 == 32'h6000;
  assign T_6821 = io_imem_resp_bits_data_0 & 32'h6018;
  assign T_6823 = T_6821 == 32'h6000;
  assign T_6825 = io_imem_resp_bits_data_0 & 32'h40003034;
  assign T_6827 = T_6825 == 32'h40000030;
  assign T_6829 = io_imem_resp_bits_data_0 & 32'h40001054;
  assign T_6831 = T_6829 == 32'h40001010;
  assign T_6834 = T_6811 | T_6815;
  assign T_6835 = T_6834 | T_6819;
  assign T_6836 = T_6835 | T_6823;
  assign T_6837 = T_6836 | T_6827;
  assign T_6838 = T_6837 | T_6831;
  assign T_6840 = io_imem_resp_bits_data_0 & 32'h2054;
  assign T_6842 = T_6840 == 32'h2010;
  assign T_6844 = io_imem_resp_bits_data_0 & 32'h40004054;
  assign T_6846 = T_6844 == 32'h4010;
  assign T_6848 = io_imem_resp_bits_data_0 & 32'h5054;
  assign T_6850 = T_6848 == 32'h4010;
  assign T_6852 = io_imem_resp_bits_data_0 & 32'h4058;
  assign T_6854 = T_6852 == 32'h4040;
  assign T_6857 = T_6842 | T_6846;
  assign T_6858 = T_6857 | T_6850;
  assign T_6859 = T_6858 | T_6854;
  assign T_6861 = io_imem_resp_bits_data_0 & 32'h6054;
  assign T_6863 = T_6861 == 32'h2010;
  assign T_6865 = io_imem_resp_bits_data_0 & 32'h40003054;
  assign T_6867 = T_6865 == 32'h40001010;
  assign T_6870 = T_6863 | T_6854;
  assign T_6871 = T_6870 | T_6827;
  assign T_6872 = T_6871 | T_6867;
  assign T_6873 = {T_6838,T_6807};
  assign T_6874 = {T_6859,T_6873};
  assign T_6875 = {T_6872,T_6874};
  assign T_6877 = io_imem_resp_bits_data_0 & 32'h605f;
  assign T_6879 = T_6877 == 32'h3;
  assign T_6881 = io_imem_resp_bits_data_0 & 32'h707f;
  assign T_6883 = T_6881 == 32'h100f;
  assign T_6886 = T_6879 | T_6564;
  assign T_6887 = T_6886 | T_6568;
  assign T_6888 = T_6887 | T_6883;
  assign T_6892 = T_6713 == 32'h20;
  assign T_6895 = T_6753 | T_6892;
  assign T_6901 = {1'h0,T_6895};
  assign T_6902 = {T_6753,T_6901};
  assign T_6903 = {1'h0,T_6902};
  assign T_6904 = {1'h0,T_6903};
  assign T_6906 = io_imem_resp_bits_data_0 & 32'h1000;
  assign T_6908 = T_6906 == 32'h1000;
  assign T_6912 = io_imem_resp_bits_data_0 & 32'h2000;
  assign T_6914 = T_6912 == 32'h2000;
  assign T_6918 = io_imem_resp_bits_data_0 & 32'h4000;
  assign T_6920 = T_6918 == 32'h4000;
  assign T_6923 = {T_6914,T_6908};
  assign T_6924 = {T_6920,T_6923};
  assign T_6930 = io_imem_resp_bits_data_0 & 32'h2000074;
  assign T_6932 = T_6930 == 32'h2000030;
  assign T_6936 = io_imem_resp_bits_data_0 & 32'h28;
  assign T_6938 = T_6936 == 32'h0;
  assign T_6940 = io_imem_resp_bits_data_0 & 32'hc;
  assign T_6942 = T_6940 == 32'h4;
  assign T_6946 = T_6709 == 32'h10;
  assign T_6948 = io_imem_resp_bits_data_0 & 32'h1010;
  assign T_6950 = T_6948 == 32'h1010;
  assign T_6952 = io_imem_resp_bits_data_0 & 32'h2010;
  assign T_6954 = T_6952 == 32'h2010;
  assign T_6957 = T_6938 | T_6942;
  assign T_6958 = T_6957 | T_6946;
  assign T_6959 = T_6958 | T_6672;
  assign T_6960 = T_6959 | T_6950;
  assign T_6961 = T_6960 | T_6954;
  assign T_6963 = io_imem_resp_bits_data_0 & 32'h1050;
  assign T_6965 = T_6963 == 32'h1050;
  assign T_6969 = io_imem_resp_bits_data_0 & 32'h2050;
  assign T_6971 = T_6969 == 32'h2050;
  assign T_6975 = io_imem_resp_bits_data_0 & 32'h3050;
  assign T_6977 = T_6975 == 32'h50;
  assign T_6980 = {T_6971,T_6965};
  assign T_6981 = {T_6977,T_6980};
  assign T_6983 = io_imem_resp_bits_data_0 & 32'h1048;
  assign T_6985 = T_6983 == 32'h1008;
  assign T_6991 = T_6983 == 32'h8;
  assign id_raddr3 = io_imem_resp_bits_data_0[31:27];
  assign id_raddr2 = io_imem_resp_bits_data_0[24:20];
  assign id_raddr1 = io_imem_resp_bits_data_0[19:15];
  assign id_waddr = io_imem_resp_bits_data_0[11:7];
  assign id_load_use = T_7744;
  assign T_6999_T_7009_addr = T_7008;
  assign T_6999_T_7009_en = 1'h1;
  `ifndef RANDOMIZE
  assign T_6999_T_7009_data = T_6999[T_6999_T_7009_addr];
  `else
  assign T_6999_T_7009_data = T_6999_T_7009_addr >= 5'h1f ? GEN_398[31:0] : T_6999[T_6999_T_7009_addr];
  `endif
  assign T_6999_T_7020_addr = T_7019;
  assign T_6999_T_7020_en = 1'h1;
  `ifndef RANDOMIZE
  assign T_6999_T_7020_data = T_6999[T_6999_T_7020_addr];
  `else
  assign T_6999_T_7020_data = T_6999_T_7020_addr >= 5'h1f ? GEN_399[31:0] : T_6999[T_6999_T_7020_addr];
  `endif
  assign T_6999_T_7648_data = rf_wdata;
  assign T_6999_T_7648_addr = T_7647;
  assign T_6999_T_7648_mask = GEN_163;
  assign T_6999_T_7648_en = GEN_163;
  assign T_7001 = GEN_166;
  assign T_7004 = id_raddr1 == 5'h0;
  assign T_7008 = ~ id_raddr1;
  assign T_7010 = T_6999_T_7009_data;
  assign T_7012 = GEN_167;
  assign T_7019 = ~ id_raddr2;
  assign T_7021 = T_6999_T_7020_data;
  assign ctrl_killd = T_7794;
  assign csr_clk = clk;
  assign csr_reset = reset;
  assign csr_io_prci_reset = io_prci_reset;
  assign csr_io_prci_id = io_prci_id;
  assign csr_io_prci_interrupts_meip = io_prci_interrupts_meip;
  assign csr_io_prci_interrupts_seip = io_prci_interrupts_seip;
  assign csr_io_prci_interrupts_debug = io_prci_interrupts_debug;
  assign csr_io_prci_interrupts_mtip = io_prci_interrupts_mtip;
  assign csr_io_prci_interrupts_msip = io_prci_interrupts_msip;
  assign csr_io_rw_addr = T_7652;
  assign csr_io_rw_cmd = T_7653;
  assign csr_io_rw_wdata = wb_reg_wdata;
  assign csr_io_exception = wb_reg_xcpt;
  assign csr_io_retire = wb_valid;
  assign csr_io_cause = wb_reg_cause;
  assign csr_io_pc = wb_reg_pc;
  assign csr_io_badaddr = T_7651;
  assign csr_io_fcsr_flags_valid = io_fpu_fcsr_flags_valid;
  assign csr_io_fcsr_flags_bits = io_fpu_fcsr_flags_bits;
  assign csr_io_rocc_cmd_ready = GEN_223;
  assign csr_io_rocc_resp_valid = GEN_224;
  assign csr_io_rocc_resp_bits_rd = GEN_225;
  assign csr_io_rocc_resp_bits_data = GEN_226;
  assign csr_io_rocc_mem_req_valid = GEN_227;
  assign csr_io_rocc_mem_req_bits_addr = GEN_228;
  assign csr_io_rocc_mem_req_bits_tag = GEN_229;
  assign csr_io_rocc_mem_req_bits_cmd = GEN_230;
  assign csr_io_rocc_mem_req_bits_typ = GEN_231;
  assign csr_io_rocc_mem_req_bits_phys = GEN_232;
  assign csr_io_rocc_mem_req_bits_data = GEN_233;
  assign csr_io_rocc_mem_s1_kill = GEN_234;
  assign csr_io_rocc_mem_s1_data = GEN_235;
  assign csr_io_rocc_mem_invalidate_lr = GEN_236;
  assign csr_io_rocc_busy = GEN_237;
  assign csr_io_rocc_interrupt = io_rocc_interrupt;
  assign csr_io_rocc_autl_acquire_valid = GEN_238;
  assign csr_io_rocc_autl_acquire_bits_addr_block = GEN_239;
  assign csr_io_rocc_autl_acquire_bits_client_xact_id = GEN_240;
  assign csr_io_rocc_autl_acquire_bits_addr_beat = GEN_241;
  assign csr_io_rocc_autl_acquire_bits_is_builtin_type = GEN_242;
  assign csr_io_rocc_autl_acquire_bits_a_type = GEN_243;
  assign csr_io_rocc_autl_acquire_bits_union = GEN_244;
  assign csr_io_rocc_autl_acquire_bits_data = GEN_245;
  assign csr_io_rocc_autl_grant_ready = GEN_246;
  assign csr_io_rocc_fpu_req_valid = GEN_247;
  assign csr_io_rocc_fpu_req_bits_cmd = GEN_248;
  assign csr_io_rocc_fpu_req_bits_ldst = GEN_249;
  assign csr_io_rocc_fpu_req_bits_wen = GEN_250;
  assign csr_io_rocc_fpu_req_bits_ren1 = GEN_251;
  assign csr_io_rocc_fpu_req_bits_ren2 = GEN_252;
  assign csr_io_rocc_fpu_req_bits_ren3 = GEN_253;
  assign csr_io_rocc_fpu_req_bits_swap12 = GEN_254;
  assign csr_io_rocc_fpu_req_bits_swap23 = GEN_255;
  assign csr_io_rocc_fpu_req_bits_single = GEN_256;
  assign csr_io_rocc_fpu_req_bits_fromint = GEN_257;
  assign csr_io_rocc_fpu_req_bits_toint = GEN_258;
  assign csr_io_rocc_fpu_req_bits_fastpipe = GEN_259;
  assign csr_io_rocc_fpu_req_bits_fma = GEN_260;
  assign csr_io_rocc_fpu_req_bits_div = GEN_261;
  assign csr_io_rocc_fpu_req_bits_sqrt = GEN_262;
  assign csr_io_rocc_fpu_req_bits_round = GEN_263;
  assign csr_io_rocc_fpu_req_bits_wflags = GEN_264;
  assign csr_io_rocc_fpu_req_bits_rm = GEN_265;
  assign csr_io_rocc_fpu_req_bits_typ = GEN_266;
  assign csr_io_rocc_fpu_req_bits_in1 = GEN_267;
  assign csr_io_rocc_fpu_req_bits_in2 = GEN_268;
  assign csr_io_rocc_fpu_req_bits_in3 = GEN_269;
  assign csr_io_rocc_fpu_resp_ready = GEN_270;
  assign id_csr_en = id_ctrl_csr != 3'h0;
  assign id_system_insn = id_ctrl_csr == 3'h4;
  assign T_7023 = id_ctrl_csr == 3'h2;
  assign T_7024 = id_ctrl_csr == 3'h3;
  assign T_7025 = T_7023 | T_7024;
  assign id_csr_ren = T_7025 & T_7004;
  assign id_csr = id_csr_ren ? 3'h5 : id_ctrl_csr;
  assign id_csr_addr = io_imem_resp_bits_data_0[31:20];
  assign T_7029 = id_csr_ren == 1'h0;
  assign T_7030 = id_csr_en & T_7029;
  assign T_7084 = id_csr_addr & 12'h46;
  assign T_7086 = T_7084 == 12'h40;
  assign T_7088 = id_csr_addr & 12'h644;
  assign T_7090 = T_7088 == 12'h240;
  assign T_7093 = T_7086 | T_7090;
  assign T_7096 = T_7093 == 1'h0;
  assign T_7097 = T_7030 & T_7096;
  assign id_csr_flush = id_system_insn | T_7097;
  assign T_7099 = id_ctrl_legal == 1'h0;
  assign T_7101 = csr_io_status_fs != 2'h0;
  assign T_7103 = T_7101 == 1'h0;
  assign T_7104 = id_ctrl_fp & T_7103;
  assign T_7105 = T_7099 | T_7104;
  assign T_7107 = csr_io_status_xs != 2'h0;
  assign T_7109 = T_7107 == 1'h0;
  assign T_7110 = id_ctrl_rocc & T_7109;
  assign id_illegal_insn = T_7105 | T_7110;
  assign id_amo_aq = io_imem_resp_bits_data_0[26];
  assign id_amo_rl = io_imem_resp_bits_data_0[25];
  assign T_7111 = id_ctrl_amo & id_amo_rl;
  assign id_fence_next = id_ctrl_fence | T_7111;
  assign T_7113 = io_dmem_ordered == 1'h0;
  assign id_mem_busy = T_7113 | io_dmem_req_valid;
  assign T_7119 = wb_reg_valid & wb_ctrl_rocc;
  assign T_7121 = id_reg_fence & id_mem_busy;
  assign T_7122 = id_fence_next | T_7121;
  assign T_7124 = id_ctrl_amo & id_amo_aq;
  assign T_7125 = T_7124 | id_ctrl_fence_i;
  assign T_7126 = id_ctrl_mem | id_ctrl_rocc;
  assign T_7127 = id_reg_fence & T_7126;
  assign T_7128 = T_7125 | T_7127;
  assign T_7129 = T_7128 | id_csr_en;
  assign T_7130 = id_mem_busy & T_7129;
  assign bpu_clk = clk;
  assign bpu_reset = reset;
  assign bpu_io_status_debug = csr_io_status_debug;
  assign bpu_io_status_prv = csr_io_status_prv;
  assign bpu_io_status_sd = csr_io_status_sd;
  assign bpu_io_status_zero3 = csr_io_status_zero3;
  assign bpu_io_status_sd_rv32 = csr_io_status_sd_rv32;
  assign bpu_io_status_zero2 = csr_io_status_zero2;
  assign bpu_io_status_vm = csr_io_status_vm;
  assign bpu_io_status_zero1 = csr_io_status_zero1;
  assign bpu_io_status_mxr = csr_io_status_mxr;
  assign bpu_io_status_pum = csr_io_status_pum;
  assign bpu_io_status_mprv = csr_io_status_mprv;
  assign bpu_io_status_xs = csr_io_status_xs;
  assign bpu_io_status_fs = csr_io_status_fs;
  assign bpu_io_status_mpp = csr_io_status_mpp;
  assign bpu_io_status_hpp = csr_io_status_hpp;
  assign bpu_io_status_spp = csr_io_status_spp;
  assign bpu_io_status_mpie = csr_io_status_mpie;
  assign bpu_io_status_hpie = csr_io_status_hpie;
  assign bpu_io_status_spie = csr_io_status_spie;
  assign bpu_io_status_upie = csr_io_status_upie;
  assign bpu_io_status_mie = csr_io_status_mie;
  assign bpu_io_status_hie = csr_io_status_hie;
  assign bpu_io_status_sie = csr_io_status_sie;
  assign bpu_io_status_uie = csr_io_status_uie;
  assign bpu_io_bp_0_control_tdrtype = csr_io_bp_0_control_tdrtype;
  assign bpu_io_bp_0_control_bpamaskmax = csr_io_bp_0_control_bpamaskmax;
  assign bpu_io_bp_0_control_reserved = csr_io_bp_0_control_reserved;
  assign bpu_io_bp_0_control_bpaction = csr_io_bp_0_control_bpaction;
  assign bpu_io_bp_0_control_bpmatch = csr_io_bp_0_control_bpmatch;
  assign bpu_io_bp_0_control_m = csr_io_bp_0_control_m;
  assign bpu_io_bp_0_control_h = csr_io_bp_0_control_h;
  assign bpu_io_bp_0_control_s = csr_io_bp_0_control_s;
  assign bpu_io_bp_0_control_u = csr_io_bp_0_control_u;
  assign bpu_io_bp_0_control_r = csr_io_bp_0_control_r;
  assign bpu_io_bp_0_control_w = csr_io_bp_0_control_w;
  assign bpu_io_bp_0_control_x = csr_io_bp_0_control_x;
  assign bpu_io_bp_0_address = csr_io_bp_0_address;
  assign bpu_io_bp_1_control_tdrtype = csr_io_bp_1_control_tdrtype;
  assign bpu_io_bp_1_control_bpamaskmax = csr_io_bp_1_control_bpamaskmax;
  assign bpu_io_bp_1_control_reserved = csr_io_bp_1_control_reserved;
  assign bpu_io_bp_1_control_bpaction = csr_io_bp_1_control_bpaction;
  assign bpu_io_bp_1_control_bpmatch = csr_io_bp_1_control_bpmatch;
  assign bpu_io_bp_1_control_m = csr_io_bp_1_control_m;
  assign bpu_io_bp_1_control_h = csr_io_bp_1_control_h;
  assign bpu_io_bp_1_control_s = csr_io_bp_1_control_s;
  assign bpu_io_bp_1_control_u = csr_io_bp_1_control_u;
  assign bpu_io_bp_1_control_r = csr_io_bp_1_control_r;
  assign bpu_io_bp_1_control_w = csr_io_bp_1_control_w;
  assign bpu_io_bp_1_control_x = csr_io_bp_1_control_x;
  assign bpu_io_bp_1_address = csr_io_bp_1_address;
  assign bpu_io_pc = io_imem_resp_bits_pc;
  assign bpu_io_ea = mem_reg_wdata;
  assign T_7134 = csr_io_interrupt | bpu_io_xcpt_if;
  assign T_7135 = T_7134 | io_imem_resp_bits_xcpt_if;
  assign id_xcpt = T_7135 | id_illegal_insn;
  assign T_7136 = io_imem_resp_bits_xcpt_if ? 2'h1 : 2'h2;
  assign T_7137 = bpu_io_xcpt_if ? 2'h3 : T_7136;
  assign id_cause = csr_io_interrupt ? csr_io_interrupt_cause : {{30'd0}, T_7137};
  assign ex_waddr = ex_reg_inst[11:7];
  assign mem_waddr = mem_reg_inst[11:7];
  assign wb_waddr = wb_reg_inst[11:7];
  assign T_7141 = ex_reg_valid & ex_ctrl_wxd;
  assign T_7142 = mem_reg_valid & mem_ctrl_wxd;
  assign T_7144 = mem_ctrl_mem == 1'h0;
  assign T_7145 = T_7142 & T_7144;
  assign T_7147 = 5'h0 == id_raddr1;
  assign T_7149 = ex_waddr == id_raddr1;
  assign T_7150 = T_7141 & T_7149;
  assign T_7151 = mem_waddr == id_raddr1;
  assign T_7152 = T_7145 & T_7151;
  assign T_7154 = T_7142 & T_7151;
  assign T_7155 = 5'h0 == id_raddr2;
  assign T_7157 = ex_waddr == id_raddr2;
  assign T_7158 = T_7141 & T_7157;
  assign T_7159 = mem_waddr == id_raddr2;
  assign T_7160 = T_7145 & T_7159;
  assign T_7162 = T_7142 & T_7159;
  assign bypass_mux_0 = 32'h0;
  assign bypass_mux_1 = mem_reg_wdata;
  assign bypass_mux_2 = wb_reg_wdata;
  assign bypass_mux_3 = io_dmem_resp_bits_data_word_bypass;
  assign T_7190 = {ex_reg_rs_msb_0,ex_reg_rs_lsb_0};
  assign GEN_0 = GEN_4;
  assign GEN_2 = 2'h1 == ex_reg_rs_lsb_0 ? bypass_mux_1 : bypass_mux_0;
  assign GEN_3 = 2'h2 == ex_reg_rs_lsb_0 ? bypass_mux_2 : GEN_2;
  assign GEN_4 = 2'h3 == ex_reg_rs_lsb_0 ? bypass_mux_3 : GEN_3;
  assign T_7191 = ex_reg_rs_bypass_0 ? GEN_0 : T_7190;
  assign T_7192 = {ex_reg_rs_msb_1,ex_reg_rs_lsb_1};
  assign GEN_1 = GEN_7;
  assign GEN_5 = 2'h1 == ex_reg_rs_lsb_1 ? bypass_mux_1 : bypass_mux_0;
  assign GEN_6 = 2'h2 == ex_reg_rs_lsb_1 ? bypass_mux_2 : GEN_5;
  assign GEN_7 = 2'h3 == ex_reg_rs_lsb_1 ? bypass_mux_3 : GEN_6;
  assign T_7193 = ex_reg_rs_bypass_1 ? GEN_1 : T_7192;
  assign T_7194 = ex_ctrl_sel_imm == 3'h5;
  assign T_7196 = ex_reg_inst[31];
  assign T_7197 = $signed(T_7196);
  assign T_7198 = T_7194 ? $signed(1'sh0) : $signed(T_7197);
  assign T_7199 = ex_ctrl_sel_imm == 3'h2;
  assign T_7200 = ex_reg_inst[30:20];
  assign T_7201 = $signed(T_7200);
  assign T_7202 = T_7199 ? $signed(T_7201) : $signed({11{T_7198}});
  assign T_7203 = ex_ctrl_sel_imm != 3'h2;
  assign T_7204 = ex_ctrl_sel_imm != 3'h3;
  assign T_7205 = T_7203 & T_7204;
  assign T_7206 = ex_reg_inst[19:12];
  assign T_7207 = $signed(T_7206);
  assign T_7208 = T_7205 ? $signed({8{T_7198}}) : $signed(T_7207);
  assign T_7211 = T_7199 | T_7194;
  assign T_7213 = ex_ctrl_sel_imm == 3'h3;
  assign T_7214 = ex_reg_inst[20];
  assign T_7215 = $signed(T_7214);
  assign T_7216 = ex_ctrl_sel_imm == 3'h1;
  assign T_7217 = ex_reg_inst[7];
  assign T_7218 = $signed(T_7217);
  assign T_7219 = T_7216 ? $signed(T_7218) : $signed(T_7198);
  assign T_7220 = T_7213 ? $signed(T_7215) : $signed(T_7219);
  assign T_7221 = T_7211 ? $signed(1'sh0) : $signed(T_7220);
  assign T_7226 = ex_reg_inst[30:25];
  assign T_7227 = T_7211 ? 6'h0 : T_7226;
  assign T_7230 = ex_ctrl_sel_imm == 3'h0;
  assign T_7232 = T_7230 | T_7216;
  assign T_7233 = ex_reg_inst[11:8];
  assign T_7235 = ex_reg_inst[19:16];
  assign T_7236 = ex_reg_inst[24:21];
  assign T_7237 = T_7194 ? T_7235 : T_7236;
  assign T_7238 = T_7232 ? T_7233 : T_7237;
  assign T_7239 = T_7199 ? 4'h0 : T_7238;
  assign T_7242 = ex_ctrl_sel_imm == 3'h4;
  assign T_7245 = ex_reg_inst[15];
  assign T_7248 = T_7194 ? T_7245 : 1'h0;
  assign T_7250 = T_7242 ? T_7214 : T_7248;
  assign T_7252 = T_7230 ? T_7217 : T_7250;
  assign T_7253 = {T_7227,T_7239};
  assign T_7254 = {T_7253,T_7252};
  assign T_7255 = $unsigned(T_7221);
  assign T_7256 = $unsigned(T_7208);
  assign T_7257 = {T_7256,T_7255};
  assign T_7258 = $unsigned(T_7202);
  assign T_7259 = $unsigned(T_7198);
  assign T_7260 = {T_7259,T_7258};
  assign T_7261 = {T_7260,T_7257};
  assign T_7262 = {T_7261,T_7254};
  assign ex_imm = $signed(T_7262);
  assign T_7264 = $signed(T_7191);
  assign T_7265 = $signed(ex_reg_pc);
  assign T_7266 = 2'h2 == ex_ctrl_sel_alu1;
  assign T_7267 = T_7266 ? $signed(T_7265) : $signed(32'sh0);
  assign T_7268 = 2'h1 == ex_ctrl_sel_alu1;
  assign ex_op1 = T_7268 ? $signed(T_7264) : $signed(T_7267);
  assign T_7270 = $signed(T_7193);
  assign T_7272 = 2'h1 == ex_ctrl_sel_alu2;
  assign T_7273 = T_7272 ? $signed(4'sh4) : $signed(4'sh0);
  assign T_7274 = 2'h3 == ex_ctrl_sel_alu2;
  assign T_7275 = T_7274 ? $signed(ex_imm) : $signed({{28{T_7273[3]}},T_7273});
  assign T_7276 = 2'h2 == ex_ctrl_sel_alu2;
  assign ex_op2 = T_7276 ? $signed(T_7270) : $signed(T_7275);
  assign alu_clk = clk;
  assign alu_reset = reset;
  assign alu_io_dw = ex_ctrl_alu_dw;
  assign alu_io_fn = ex_ctrl_alu_fn;
  assign alu_io_in2 = T_7277;
  assign alu_io_in1 = T_7278;
  assign T_7277 = $unsigned(ex_op2);
  assign T_7278 = $unsigned(ex_op1);
  assign div_clk = clk;
  assign div_reset = reset;
  assign div_io_req_valid = T_7279;
  assign div_io_req_bits_fn = ex_ctrl_alu_fn;
  assign div_io_req_bits_dw = ex_ctrl_alu_dw;
  assign div_io_req_bits_in1 = T_7191;
  assign div_io_req_bits_in2 = T_7193;
  assign div_io_req_bits_tag = ex_waddr;
  assign div_io_kill = T_7599;
  assign div_io_resp_ready = GEN_149;
  assign T_7279 = ex_reg_valid & ex_ctrl_div;
  assign T_7281 = ctrl_killd == 1'h0;
  assign T_7283 = take_pc_mem_wb == 1'h0;
  assign T_7284 = T_7283 & io_imem_resp_valid;
  assign T_7285 = T_7284 & io_imem_resp_bits_replay;
  assign T_7288 = T_7281 & id_xcpt;
  assign T_7292 = T_7284 & csr_io_interrupt;
  assign GEN_8 = id_xcpt ? id_cause : ex_reg_cause;
  assign GEN_9 = io_imem_btb_resp_valid ? io_imem_btb_resp_bits_taken : ex_reg_btb_resp_taken;
  assign GEN_10 = io_imem_btb_resp_valid ? io_imem_btb_resp_bits_mask : ex_reg_btb_resp_mask;
  assign GEN_11 = io_imem_btb_resp_valid ? io_imem_btb_resp_bits_bridx : ex_reg_btb_resp_bridx;
  assign GEN_12 = io_imem_btb_resp_valid ? io_imem_btb_resp_bits_target : ex_reg_btb_resp_target;
  assign GEN_13 = io_imem_btb_resp_valid ? io_imem_btb_resp_bits_entry : ex_reg_btb_resp_entry;
  assign GEN_14 = io_imem_btb_resp_valid ? io_imem_btb_resp_bits_bht_history : ex_reg_btb_resp_bht_history;
  assign GEN_15 = io_imem_btb_resp_valid ? io_imem_btb_resp_bits_bht_value : ex_reg_btb_resp_bht_value;
  assign T_7295 = id_ctrl_fence_i | id_csr_flush;
  assign T_7296 = T_7295 | csr_io_singleStep;
  assign T_7297 = id_ctrl_jalr & csr_io_status_debug;
  assign GEN_16 = T_7297 ? 1'h1 : T_7296;
  assign GEN_17 = T_7297 ? 1'h1 : id_ctrl_fence_i;
  assign T_7300 = T_7147 | T_7150;
  assign T_7301 = T_7300 | T_7152;
  assign T_7302 = T_7301 | T_7154;
  assign T_7307 = T_7152 ? 2'h2 : 2'h3;
  assign T_7308 = T_7150 ? 2'h1 : T_7307;
  assign T_7309 = T_7147 ? 2'h0 : T_7308;
  assign T_7311 = T_7302 == 1'h0;
  assign T_7312 = id_ctrl_rxs1 & T_7311;
  assign T_7313 = T_7001[1:0];
  assign T_7314 = T_7001[31:2];
  assign GEN_18 = T_7312 ? T_7313 : T_7309;
  assign GEN_19 = T_7312 ? T_7314 : ex_reg_rs_msb_0;
  assign T_7315 = T_7155 | T_7158;
  assign T_7316 = T_7315 | T_7160;
  assign T_7317 = T_7316 | T_7162;
  assign T_7322 = T_7160 ? 2'h2 : 2'h3;
  assign T_7323 = T_7158 ? 2'h1 : T_7322;
  assign T_7324 = T_7155 ? 2'h0 : T_7323;
  assign T_7326 = T_7317 == 1'h0;
  assign T_7327 = id_ctrl_rxs2 & T_7326;
  assign T_7328 = T_7012[1:0];
  assign T_7329 = T_7012[31:2];
  assign GEN_20 = T_7327 ? T_7328 : T_7324;
  assign GEN_21 = T_7327 ? T_7329 : ex_reg_rs_msb_1;
  assign GEN_22 = T_7281 ? id_ctrl_legal : ex_ctrl_legal;
  assign GEN_23 = T_7281 ? id_ctrl_fp : ex_ctrl_fp;
  assign GEN_24 = T_7281 ? id_ctrl_rocc : ex_ctrl_rocc;
  assign GEN_25 = T_7281 ? id_ctrl_branch : ex_ctrl_branch;
  assign GEN_26 = T_7281 ? id_ctrl_jal : ex_ctrl_jal;
  assign GEN_27 = T_7281 ? id_ctrl_jalr : ex_ctrl_jalr;
  assign GEN_28 = T_7281 ? id_ctrl_rxs2 : ex_ctrl_rxs2;
  assign GEN_29 = T_7281 ? id_ctrl_rxs1 : ex_ctrl_rxs1;
  assign GEN_30 = T_7281 ? id_ctrl_sel_alu2 : ex_ctrl_sel_alu2;
  assign GEN_31 = T_7281 ? id_ctrl_sel_alu1 : ex_ctrl_sel_alu1;
  assign GEN_32 = T_7281 ? id_ctrl_sel_imm : ex_ctrl_sel_imm;
  assign GEN_33 = T_7281 ? id_ctrl_alu_dw : ex_ctrl_alu_dw;
  assign GEN_34 = T_7281 ? id_ctrl_alu_fn : ex_ctrl_alu_fn;
  assign GEN_35 = T_7281 ? id_ctrl_mem : ex_ctrl_mem;
  assign GEN_36 = T_7281 ? id_ctrl_mem_cmd : ex_ctrl_mem_cmd;
  assign GEN_37 = T_7281 ? id_ctrl_mem_type : ex_ctrl_mem_type;
  assign GEN_38 = T_7281 ? id_ctrl_rfs1 : ex_ctrl_rfs1;
  assign GEN_39 = T_7281 ? id_ctrl_rfs2 : ex_ctrl_rfs2;
  assign GEN_40 = T_7281 ? id_ctrl_rfs3 : ex_ctrl_rfs3;
  assign GEN_41 = T_7281 ? id_ctrl_wfd : ex_ctrl_wfd;
  assign GEN_42 = T_7281 ? id_ctrl_div : ex_ctrl_div;
  assign GEN_43 = T_7281 ? id_ctrl_wxd : ex_ctrl_wxd;
  assign GEN_44 = T_7281 ? id_csr : ex_ctrl_csr;
  assign GEN_45 = T_7281 ? GEN_17 : ex_ctrl_fence_i;
  assign GEN_46 = T_7281 ? id_ctrl_fence : ex_ctrl_fence;
  assign GEN_47 = T_7281 ? id_ctrl_amo : ex_ctrl_amo;
  assign GEN_48 = T_7281 ? io_imem_btb_resp_valid : ex_reg_btb_hit;
  assign GEN_49 = T_7281 ? GEN_9 : ex_reg_btb_resp_taken;
  assign GEN_50 = T_7281 ? GEN_10 : ex_reg_btb_resp_mask;
  assign GEN_51 = T_7281 ? GEN_11 : ex_reg_btb_resp_bridx;
  assign GEN_52 = T_7281 ? GEN_12 : ex_reg_btb_resp_target;
  assign GEN_53 = T_7281 ? GEN_13 : ex_reg_btb_resp_entry;
  assign GEN_54 = T_7281 ? GEN_14 : ex_reg_btb_resp_bht_history;
  assign GEN_55 = T_7281 ? GEN_15 : ex_reg_btb_resp_bht_value;
  assign GEN_56 = T_7281 ? GEN_16 : ex_reg_flush_pipe;
  assign GEN_57 = T_7281 ? id_load_use : ex_reg_load_use;
  assign GEN_58 = T_7281 ? T_7302 : ex_reg_rs_bypass_0;
  assign GEN_59 = T_7281 ? GEN_18 : ex_reg_rs_lsb_0;
  assign GEN_60 = T_7281 ? GEN_19 : ex_reg_rs_msb_0;
  assign GEN_61 = T_7281 ? T_7317 : ex_reg_rs_bypass_1;
  assign GEN_62 = T_7281 ? GEN_20 : ex_reg_rs_lsb_1;
  assign GEN_63 = T_7281 ? GEN_21 : ex_reg_rs_msb_1;
  assign T_7332 = T_7281 | csr_io_interrupt;
  assign T_7333 = T_7332 | io_imem_resp_bits_replay;
  assign GEN_64 = T_7333 ? io_imem_resp_bits_data_0 : ex_reg_inst;
  assign GEN_65 = T_7333 ? io_imem_resp_bits_pc : ex_reg_pc;
  assign T_7334 = ex_reg_valid | ex_reg_replay;
  assign ex_pc_valid = T_7334 | ex_reg_xcpt_interrupt;
  assign T_7336 = io_dmem_resp_valid == 1'h0;
  assign wb_dcache_miss = wb_ctrl_mem & T_7336;
  assign T_7338 = io_dmem_req_ready == 1'h0;
  assign T_7339 = ex_ctrl_mem & T_7338;
  assign T_7341 = div_io_req_ready == 1'h0;
  assign T_7342 = ex_ctrl_div & T_7341;
  assign replay_ex_structural = T_7339 | T_7342;
  assign replay_ex_load_use = wb_dcache_miss & ex_reg_load_use;
  assign T_7343 = replay_ex_structural | replay_ex_load_use;
  assign T_7344 = ex_reg_valid & T_7343;
  assign replay_ex = ex_reg_replay | T_7344;
  assign T_7345 = take_pc_mem_wb | replay_ex;
  assign T_7347 = ex_reg_valid == 1'h0;
  assign ctrl_killx = T_7345 | T_7347;
  assign T_7348 = ex_ctrl_mem_cmd == 5'h7;
  assign T_7354_0 = 3'h0;
  assign T_7354_1 = 3'h4;
  assign T_7354_2 = 3'h1;
  assign T_7354_3 = 3'h5;
  assign T_7356 = T_7354_0 == ex_ctrl_mem_type;
  assign T_7357 = T_7354_1 == ex_ctrl_mem_type;
  assign T_7358 = T_7354_2 == ex_ctrl_mem_type;
  assign T_7359 = T_7354_3 == ex_ctrl_mem_type;
  assign T_7362 = T_7356 | T_7357;
  assign T_7363 = T_7362 | T_7358;
  assign T_7364 = T_7363 | T_7359;
  assign ex_slow_bypass = T_7348 | T_7364;
  assign T_7365 = ex_reg_xcpt_interrupt | ex_reg_xcpt;
  assign T_7366 = ex_ctrl_fp & io_fpu_illegal_rm;
  assign ex_xcpt = T_7365 | T_7366;
  assign ex_cause = T_7365 ? ex_reg_cause : 32'h2;
  assign mem_br_taken = mem_reg_wdata[0];
  assign T_7368 = $signed(mem_reg_pc);
  assign T_7369 = mem_ctrl_branch & mem_br_taken;
  assign T_7372 = mem_reg_inst[31];
  assign T_7373 = $signed(T_7372);
  assign T_7378 = {11{T_7373}};
  assign T_7382 = mem_reg_inst[19:12];
  assign T_7383 = $signed(T_7382);
  assign T_7384 = {8{T_7373}};
  assign T_7390 = mem_reg_inst[20];
  assign T_7391 = $signed(T_7390);
  assign T_7393 = mem_reg_inst[7];
  assign T_7394 = $signed(T_7393);
  assign T_7402 = mem_reg_inst[30:25];
  assign T_7409 = mem_reg_inst[11:8];
  assign T_7412 = mem_reg_inst[24:21];
  assign T_7429 = {T_7402,T_7409};
  assign T_7430 = {T_7429,1'h0};
  assign T_7431 = $unsigned(T_7394);
  assign T_7432 = $unsigned(T_7384);
  assign T_7433 = {T_7432,T_7431};
  assign T_7434 = $unsigned(T_7378);
  assign T_7435 = $unsigned(T_7373);
  assign T_7436 = {T_7435,T_7434};
  assign T_7437 = {T_7436,T_7433};
  assign T_7438 = {T_7437,T_7430};
  assign T_7439 = $signed(T_7438);
  assign T_7499 = {T_7402,T_7412};
  assign T_7500 = {T_7499,1'h0};
  assign T_7501 = $unsigned(T_7391);
  assign T_7502 = $unsigned(T_7383);
  assign T_7503 = {T_7502,T_7501};
  assign T_7507 = {T_7436,T_7503};
  assign T_7508 = {T_7507,T_7500};
  assign T_7509 = $signed(T_7508);
  assign T_7511 = mem_ctrl_jal ? $signed(T_7509) : $signed(32'sh4);
  assign T_7512 = T_7369 ? $signed(T_7439) : $signed(T_7511);
  assign T_7513 = $signed(T_7368) + $signed(T_7512);
  assign T_7514 = T_7513[31:0];
  assign mem_br_target = $signed(T_7514);
  assign T_7515 = $signed(mem_reg_wdata);
  assign T_7516 = mem_ctrl_jalr ? $signed(mem_br_target) : $signed(T_7515);
  assign mem_int_wdata = $unsigned(T_7516);
  assign T_7518 = mem_ctrl_jalr ? $signed(T_7515) : $signed(mem_br_target);
  assign T_7520 = $signed(T_7518) & $signed(32'shfffffffe);
  assign T_7521 = $signed(T_7520);
  assign mem_npc = $unsigned(T_7521);
  assign T_7522 = mem_npc != ex_reg_pc;
  assign T_7523 = mem_npc != io_imem_resp_bits_pc;
  assign T_7525 = io_imem_resp_valid ? T_7523 : 1'h1;
  assign mem_wrong_npc = ex_pc_valid ? T_7522 : T_7525;
  assign mem_npc_misaligned = mem_npc[1];
  assign T_7528 = T_7369 | mem_ctrl_jalr;
  assign mem_misprediction = T_7528 | mem_ctrl_jal;
  assign T_7529 = mem_misprediction | mem_reg_flush_pipe;
  assign want_take_pc_mem = mem_reg_valid & T_7529;
  assign T_7531 = mem_npc_misaligned == 1'h0;
  assign T_7532 = want_take_pc_mem & T_7531;
  assign T_7534 = ctrl_killx == 1'h0;
  assign T_7537 = T_7283 & replay_ex;
  assign T_7540 = T_7534 & ex_xcpt;
  assign T_7543 = T_7283 & ex_reg_xcpt_interrupt;
  assign GEN_66 = ex_xcpt ? ex_cause : mem_reg_cause;
  assign T_7544 = ex_ctrl_mem_cmd == 5'h0;
  assign T_7545 = ex_ctrl_mem_cmd == 5'h6;
  assign T_7546 = T_7544 | T_7545;
  assign T_7548 = T_7546 | T_7348;
  assign T_7549 = ex_ctrl_mem_cmd[3];
  assign T_7550 = ex_ctrl_mem_cmd == 5'h4;
  assign T_7551 = T_7549 | T_7550;
  assign T_7552 = T_7548 | T_7551;
  assign T_7553 = ex_ctrl_mem & T_7552;
  assign T_7554 = ex_ctrl_mem_cmd == 5'h1;
  assign T_7556 = T_7554 | T_7348;
  assign T_7560 = T_7556 | T_7551;
  assign T_7561 = ex_ctrl_mem & T_7560;
  assign GEN_67 = ex_reg_btb_hit ? ex_reg_btb_resp_taken : mem_reg_btb_resp_taken;
  assign GEN_68 = ex_reg_btb_hit ? ex_reg_btb_resp_mask : mem_reg_btb_resp_mask;
  assign GEN_69 = ex_reg_btb_hit ? ex_reg_btb_resp_bridx : mem_reg_btb_resp_bridx;
  assign GEN_70 = ex_reg_btb_hit ? ex_reg_btb_resp_target : mem_reg_btb_resp_target;
  assign GEN_71 = ex_reg_btb_hit ? ex_reg_btb_resp_entry : mem_reg_btb_resp_entry;
  assign GEN_72 = ex_reg_btb_hit ? ex_reg_btb_resp_bht_history : mem_reg_btb_resp_bht_history;
  assign GEN_73 = ex_reg_btb_hit ? ex_reg_btb_resp_bht_value : mem_reg_btb_resp_bht_value;
  assign T_7562 = ex_ctrl_mem | ex_ctrl_rocc;
  assign T_7563 = ex_ctrl_rxs2 & T_7562;
  assign GEN_74 = T_7563 ? T_7193 : mem_reg_rs2;
  assign GEN_75 = ex_pc_valid ? ex_ctrl_legal : mem_ctrl_legal;
  assign GEN_76 = ex_pc_valid ? ex_ctrl_fp : mem_ctrl_fp;
  assign GEN_77 = ex_pc_valid ? ex_ctrl_rocc : mem_ctrl_rocc;
  assign GEN_78 = ex_pc_valid ? ex_ctrl_branch : mem_ctrl_branch;
  assign GEN_79 = ex_pc_valid ? ex_ctrl_jal : mem_ctrl_jal;
  assign GEN_80 = ex_pc_valid ? ex_ctrl_jalr : mem_ctrl_jalr;
  assign GEN_81 = ex_pc_valid ? ex_ctrl_rxs2 : mem_ctrl_rxs2;
  assign GEN_82 = ex_pc_valid ? ex_ctrl_rxs1 : mem_ctrl_rxs1;
  assign GEN_83 = ex_pc_valid ? ex_ctrl_sel_alu2 : mem_ctrl_sel_alu2;
  assign GEN_84 = ex_pc_valid ? ex_ctrl_sel_alu1 : mem_ctrl_sel_alu1;
  assign GEN_85 = ex_pc_valid ? ex_ctrl_sel_imm : mem_ctrl_sel_imm;
  assign GEN_86 = ex_pc_valid ? ex_ctrl_alu_dw : mem_ctrl_alu_dw;
  assign GEN_87 = ex_pc_valid ? ex_ctrl_alu_fn : mem_ctrl_alu_fn;
  assign GEN_88 = ex_pc_valid ? ex_ctrl_mem : mem_ctrl_mem;
  assign GEN_89 = ex_pc_valid ? ex_ctrl_mem_cmd : mem_ctrl_mem_cmd;
  assign GEN_90 = ex_pc_valid ? ex_ctrl_mem_type : mem_ctrl_mem_type;
  assign GEN_91 = ex_pc_valid ? ex_ctrl_rfs1 : mem_ctrl_rfs1;
  assign GEN_92 = ex_pc_valid ? ex_ctrl_rfs2 : mem_ctrl_rfs2;
  assign GEN_93 = ex_pc_valid ? ex_ctrl_rfs3 : mem_ctrl_rfs3;
  assign GEN_94 = ex_pc_valid ? ex_ctrl_wfd : mem_ctrl_wfd;
  assign GEN_95 = ex_pc_valid ? ex_ctrl_div : mem_ctrl_div;
  assign GEN_96 = ex_pc_valid ? ex_ctrl_wxd : mem_ctrl_wxd;
  assign GEN_97 = ex_pc_valid ? ex_ctrl_csr : mem_ctrl_csr;
  assign GEN_98 = ex_pc_valid ? ex_ctrl_fence_i : mem_ctrl_fence_i;
  assign GEN_99 = ex_pc_valid ? ex_ctrl_fence : mem_ctrl_fence;
  assign GEN_100 = ex_pc_valid ? ex_ctrl_amo : mem_ctrl_amo;
  assign GEN_101 = ex_pc_valid ? T_7553 : mem_reg_load;
  assign GEN_102 = ex_pc_valid ? T_7561 : mem_reg_store;
  assign GEN_103 = ex_pc_valid ? ex_reg_btb_hit : mem_reg_btb_hit;
  assign GEN_104 = ex_pc_valid ? GEN_67 : mem_reg_btb_resp_taken;
  assign GEN_105 = ex_pc_valid ? GEN_68 : mem_reg_btb_resp_mask;
  assign GEN_106 = ex_pc_valid ? GEN_69 : mem_reg_btb_resp_bridx;
  assign GEN_107 = ex_pc_valid ? GEN_70 : mem_reg_btb_resp_target;
  assign GEN_108 = ex_pc_valid ? GEN_71 : mem_reg_btb_resp_entry;
  assign GEN_109 = ex_pc_valid ? GEN_72 : mem_reg_btb_resp_bht_history;
  assign GEN_110 = ex_pc_valid ? GEN_73 : mem_reg_btb_resp_bht_value;
  assign GEN_111 = ex_pc_valid ? ex_reg_flush_pipe : mem_reg_flush_pipe;
  assign GEN_112 = ex_pc_valid ? ex_slow_bypass : mem_reg_slow_bypass;
  assign GEN_113 = ex_pc_valid ? ex_reg_inst : mem_reg_inst;
  assign GEN_114 = ex_pc_valid ? ex_reg_pc : mem_reg_pc;
  assign GEN_115 = ex_pc_valid ? alu_io_out : mem_reg_wdata;
  assign GEN_116 = ex_pc_valid ? GEN_74 : mem_reg_rs2;
  assign T_7564 = mem_reg_load & bpu_io_xcpt_ld;
  assign T_7566 = mem_reg_store & bpu_io_xcpt_st;
  assign T_7568 = want_take_pc_mem & mem_npc_misaligned;
  assign T_7570 = mem_ctrl_mem & io_dmem_xcpt_ma_st;
  assign T_7572 = mem_ctrl_mem & io_dmem_xcpt_ma_ld;
  assign T_7574 = mem_ctrl_mem & io_dmem_xcpt_pf_st;
  assign T_7576 = mem_ctrl_mem & io_dmem_xcpt_pf_ld;
  assign T_7578 = T_7564 | T_7566;
  assign T_7579 = T_7578 | T_7568;
  assign T_7580 = T_7579 | T_7570;
  assign T_7581 = T_7580 | T_7572;
  assign T_7582 = T_7581 | T_7574;
  assign mem_new_xcpt = T_7582 | T_7576;
  assign T_7583 = T_7574 ? 3'h7 : 3'h5;
  assign T_7584 = T_7572 ? 3'h4 : T_7583;
  assign T_7585 = T_7570 ? 3'h6 : T_7584;
  assign T_7586 = T_7568 ? 3'h0 : T_7585;
  assign T_7587 = T_7566 ? 3'h3 : T_7586;
  assign mem_new_cause = T_7564 ? 3'h3 : T_7587;
  assign T_7588 = mem_reg_xcpt_interrupt | mem_reg_xcpt;
  assign T_7589 = mem_reg_valid & mem_new_xcpt;
  assign mem_xcpt = T_7588 | T_7589;
  assign mem_cause = T_7588 ? mem_reg_cause : {{29'd0}, mem_new_cause};
  assign dcache_kill_mem = T_7142 & io_dmem_replay_next;
  assign T_7591 = mem_reg_valid & mem_ctrl_fp;
  assign fpu_kill_mem = T_7591 & io_fpu_nack_mem;
  assign T_7592 = dcache_kill_mem | mem_reg_replay;
  assign replay_mem = T_7592 | fpu_kill_mem;
  assign T_7593 = dcache_kill_mem | take_pc_wb;
  assign T_7594 = T_7593 | mem_reg_xcpt;
  assign T_7596 = mem_reg_valid == 1'h0;
  assign killm_common = T_7594 | T_7596;
  assign T_7597 = div_io_req_ready & div_io_req_valid;
  assign T_7599 = killm_common & T_7598;
  assign T_7600 = killm_common | mem_xcpt;
  assign ctrl_killm = T_7600 | fpu_kill_mem;
  assign T_7602 = ctrl_killm == 1'h0;
  assign T_7604 = take_pc_wb == 1'h0;
  assign T_7605 = replay_mem & T_7604;
  assign T_7608 = mem_xcpt & T_7604;
  assign T_7612 = T_7588 == 1'h0;
  assign T_7613 = T_7589 & T_7612;
  assign GEN_117 = mem_xcpt ? mem_cause : wb_reg_cause;
  assign T_7614 = mem_reg_valid | mem_reg_replay;
  assign T_7615 = T_7614 | mem_reg_xcpt_interrupt;
  assign T_7616 = mem_ctrl_fp & mem_ctrl_wxd;
  assign T_7617 = T_7616 ? io_fpu_toint_data : mem_int_wdata;
  assign GEN_118 = mem_ctrl_rocc ? mem_reg_rs2 : wb_reg_rs2;
  assign GEN_119 = T_7615 ? mem_ctrl_legal : wb_ctrl_legal;
  assign GEN_120 = T_7615 ? mem_ctrl_fp : wb_ctrl_fp;
  assign GEN_121 = T_7615 ? mem_ctrl_rocc : wb_ctrl_rocc;
  assign GEN_122 = T_7615 ? mem_ctrl_branch : wb_ctrl_branch;
  assign GEN_123 = T_7615 ? mem_ctrl_jal : wb_ctrl_jal;
  assign GEN_124 = T_7615 ? mem_ctrl_jalr : wb_ctrl_jalr;
  assign GEN_125 = T_7615 ? mem_ctrl_rxs2 : wb_ctrl_rxs2;
  assign GEN_126 = T_7615 ? mem_ctrl_rxs1 : wb_ctrl_rxs1;
  assign GEN_127 = T_7615 ? mem_ctrl_sel_alu2 : wb_ctrl_sel_alu2;
  assign GEN_128 = T_7615 ? mem_ctrl_sel_alu1 : wb_ctrl_sel_alu1;
  assign GEN_129 = T_7615 ? mem_ctrl_sel_imm : wb_ctrl_sel_imm;
  assign GEN_130 = T_7615 ? mem_ctrl_alu_dw : wb_ctrl_alu_dw;
  assign GEN_131 = T_7615 ? mem_ctrl_alu_fn : wb_ctrl_alu_fn;
  assign GEN_132 = T_7615 ? mem_ctrl_mem : wb_ctrl_mem;
  assign GEN_133 = T_7615 ? mem_ctrl_mem_cmd : wb_ctrl_mem_cmd;
  assign GEN_134 = T_7615 ? mem_ctrl_mem_type : wb_ctrl_mem_type;
  assign GEN_135 = T_7615 ? mem_ctrl_rfs1 : wb_ctrl_rfs1;
  assign GEN_136 = T_7615 ? mem_ctrl_rfs2 : wb_ctrl_rfs2;
  assign GEN_137 = T_7615 ? mem_ctrl_rfs3 : wb_ctrl_rfs3;
  assign GEN_138 = T_7615 ? mem_ctrl_wfd : wb_ctrl_wfd;
  assign GEN_139 = T_7615 ? mem_ctrl_div : wb_ctrl_div;
  assign GEN_140 = T_7615 ? mem_ctrl_wxd : wb_ctrl_wxd;
  assign GEN_141 = T_7615 ? mem_ctrl_csr : wb_ctrl_csr;
  assign GEN_142 = T_7615 ? mem_ctrl_fence_i : wb_ctrl_fence_i;
  assign GEN_143 = T_7615 ? mem_ctrl_fence : wb_ctrl_fence;
  assign GEN_144 = T_7615 ? mem_ctrl_amo : wb_ctrl_amo;
  assign GEN_145 = T_7615 ? T_7617 : wb_reg_wdata;
  assign GEN_146 = T_7615 ? GEN_118 : wb_reg_rs2;
  assign GEN_147 = T_7615 ? mem_reg_inst : wb_reg_inst;
  assign GEN_148 = T_7615 ? mem_reg_pc : wb_reg_pc;
  assign T_7618 = wb_ctrl_div | wb_dcache_miss;
  assign wb_set_sboard = T_7618 | wb_ctrl_rocc;
  assign replay_wb_common = io_dmem_s2_nack | wb_reg_replay;
  assign T_7621 = io_rocc_cmd_ready == 1'h0;
  assign replay_wb_rocc = T_7119 & T_7621;
  assign replay_wb = replay_wb_common | replay_wb_rocc;
  assign wb_xcpt = wb_reg_xcpt | csr_io_csr_xcpt;
  assign T_7622 = replay_wb | wb_xcpt;
  assign T_7623 = T_7622 | csr_io_eret;
  assign T_7624 = io_dmem_resp_bits_tag[0];
  assign dmem_resp_xpu = T_7624 == 1'h0;
  assign dmem_resp_waddr = io_dmem_resp_bits_tag[8:1];
  assign dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data;
  assign dmem_resp_replay = dmem_resp_valid & io_dmem_resp_bits_replay;
  assign T_7628 = wb_reg_valid & wb_ctrl_wxd;
  assign T_7630 = T_7628 == 1'h0;
  assign ll_wdata = div_io_resp_bits_data;
  assign ll_waddr = GEN_150;
  assign T_7631 = div_io_resp_ready & div_io_resp_valid;
  assign ll_wen = GEN_151;
  assign T_7632 = dmem_resp_replay & dmem_resp_xpu;
  assign GEN_149 = T_7632 ? 1'h0 : T_7630;
  assign GEN_150 = T_7632 ? dmem_resp_waddr : {{3'd0}, div_io_resp_bits_tag};
  assign GEN_151 = T_7632 ? 1'h1 : T_7631;
  assign T_7636 = replay_wb == 1'h0;
  assign T_7637 = wb_reg_valid & T_7636;
  assign T_7639 = wb_xcpt == 1'h0;
  assign wb_valid = T_7637 & T_7639;
  assign wb_wen = wb_valid & wb_ctrl_wxd;
  assign rf_wen = wb_wen | ll_wen;
  assign rf_waddr = ll_wen ? ll_waddr : {{3'd0}, wb_waddr};
  assign T_7640 = dmem_resp_valid & dmem_resp_xpu;
  assign T_7641 = wb_ctrl_csr != 3'h0;
  assign T_7642 = T_7641 ? csr_io_rw_rdata : wb_reg_wdata;
  assign T_7643 = ll_wen ? ll_wdata : T_7642;
  assign rf_wdata = T_7640 ? io_dmem_resp_bits_data : T_7643;
  assign T_7645 = rf_waddr != 8'h0;
  assign T_7646 = rf_waddr[4:0];
  assign T_7647 = ~ T_7646;
  assign GEN_170 = {{3'd0}, id_raddr1};
  assign T_7649 = rf_waddr == GEN_170;
  assign GEN_152 = T_7649 ? rf_wdata : T_7010;
  assign GEN_171 = {{3'd0}, id_raddr2};
  assign T_7650 = rf_waddr == GEN_171;
  assign GEN_153 = T_7650 ? rf_wdata : T_7021;
  assign GEN_159 = T_7645 ? GEN_152 : T_7010;
  assign GEN_160 = T_7645 ? GEN_153 : T_7021;
  assign GEN_163 = rf_wen ? T_7645 : 1'h0;
  assign GEN_166 = rf_wen ? GEN_159 : T_7010;
  assign GEN_167 = rf_wen ? GEN_160 : T_7021;
  assign T_7651 = wb_reg_mem_xcpt ? wb_reg_wdata : wb_reg_pc;
  assign T_7652 = wb_reg_inst[31:20];
  assign T_7653 = wb_reg_valid ? wb_ctrl_csr : 3'h0;
  assign T_7655 = id_raddr1 != 5'h0;
  assign T_7656 = id_ctrl_rxs1 & T_7655;
  assign T_7658 = id_raddr2 != 5'h0;
  assign T_7659 = id_ctrl_rxs2 & T_7658;
  assign T_7661 = id_waddr != 5'h0;
  assign T_7662 = id_ctrl_wxd & T_7661;
  assign T_7667 = 256'h1 << ll_waddr;
  assign T_7669 = ll_wen ? T_7667 : 256'h0;
  assign T_7670 = ~ T_7669;
  assign GEN_172 = {{224'd0}, T_7664};
  assign T_7671 = GEN_172 & T_7670;
  assign GEN_168 = ll_wen ? T_7671 : {{224'd0}, T_7664};
  assign T_7673 = T_7664 >> id_raddr1;
  assign T_7674 = T_7673[0];
  assign T_7675 = T_7656 & T_7674;
  assign T_7676 = T_7664 >> id_raddr2;
  assign T_7677 = T_7676[0];
  assign T_7678 = T_7659 & T_7677;
  assign T_7679 = T_7664 >> id_waddr;
  assign T_7680 = T_7679[0];
  assign T_7681 = T_7662 & T_7680;
  assign T_7682 = T_7675 | T_7678;
  assign id_sboard_hazard = T_7682 | T_7681;
  assign T_7683 = wb_set_sboard & wb_wen;
  assign T_7685 = 32'h1 << wb_waddr;
  assign T_7687 = T_7683 ? T_7685 : 32'h0;
  assign GEN_173 = {{224'd0}, T_7687};
  assign T_7688 = T_7671 | GEN_173;
  assign T_7689 = ll_wen | T_7683;
  assign GEN_169 = T_7689 ? T_7688 : GEN_168;
  assign T_7690 = ex_ctrl_csr != 3'h0;
  assign T_7691 = T_7690 | ex_ctrl_jalr;
  assign T_7692 = T_7691 | ex_ctrl_mem;
  assign T_7693 = T_7692 | ex_ctrl_div;
  assign T_7694 = T_7693 | ex_ctrl_fp;
  assign ex_cannot_bypass = T_7694 | ex_ctrl_rocc;
  assign T_7695 = id_raddr1 == ex_waddr;
  assign T_7696 = T_7656 & T_7695;
  assign T_7697 = id_raddr2 == ex_waddr;
  assign T_7698 = T_7659 & T_7697;
  assign T_7699 = id_waddr == ex_waddr;
  assign T_7700 = T_7662 & T_7699;
  assign T_7701 = T_7696 | T_7698;
  assign T_7702 = T_7701 | T_7700;
  assign data_hazard_ex = ex_ctrl_wxd & T_7702;
  assign T_7704 = io_fpu_dec_ren1 & T_7695;
  assign T_7706 = io_fpu_dec_ren2 & T_7697;
  assign T_7707 = id_raddr3 == ex_waddr;
  assign T_7708 = io_fpu_dec_ren3 & T_7707;
  assign T_7710 = io_fpu_dec_wen & T_7699;
  assign T_7711 = T_7704 | T_7706;
  assign T_7712 = T_7711 | T_7708;
  assign T_7713 = T_7712 | T_7710;
  assign fp_data_hazard_ex = ex_ctrl_wfd & T_7713;
  assign T_7714 = data_hazard_ex & ex_cannot_bypass;
  assign T_7715 = T_7714 | fp_data_hazard_ex;
  assign id_ex_hazard = ex_reg_valid & T_7715;
  assign T_7717 = mem_ctrl_csr != 3'h0;
  assign T_7718 = mem_ctrl_mem & mem_reg_slow_bypass;
  assign T_7719 = T_7717 | T_7718;
  assign T_7720 = T_7719 | mem_ctrl_div;
  assign T_7721 = T_7720 | mem_ctrl_fp;
  assign mem_cannot_bypass = T_7721 | mem_ctrl_rocc;
  assign T_7722 = id_raddr1 == mem_waddr;
  assign T_7723 = T_7656 & T_7722;
  assign T_7724 = id_raddr2 == mem_waddr;
  assign T_7725 = T_7659 & T_7724;
  assign T_7726 = id_waddr == mem_waddr;
  assign T_7727 = T_7662 & T_7726;
  assign T_7728 = T_7723 | T_7725;
  assign T_7729 = T_7728 | T_7727;
  assign data_hazard_mem = mem_ctrl_wxd & T_7729;
  assign T_7731 = io_fpu_dec_ren1 & T_7722;
  assign T_7733 = io_fpu_dec_ren2 & T_7724;
  assign T_7734 = id_raddr3 == mem_waddr;
  assign T_7735 = io_fpu_dec_ren3 & T_7734;
  assign T_7737 = io_fpu_dec_wen & T_7726;
  assign T_7738 = T_7731 | T_7733;
  assign T_7739 = T_7738 | T_7735;
  assign T_7740 = T_7739 | T_7737;
  assign fp_data_hazard_mem = mem_ctrl_wfd & T_7740;
  assign T_7741 = data_hazard_mem & mem_cannot_bypass;
  assign T_7742 = T_7741 | fp_data_hazard_mem;
  assign id_mem_hazard = mem_reg_valid & T_7742;
  assign T_7743 = mem_reg_valid & data_hazard_mem;
  assign T_7744 = T_7743 & mem_ctrl_mem;
  assign T_7745 = id_raddr1 == wb_waddr;
  assign T_7746 = T_7656 & T_7745;
  assign T_7747 = id_raddr2 == wb_waddr;
  assign T_7748 = T_7659 & T_7747;
  assign T_7749 = id_waddr == wb_waddr;
  assign T_7750 = T_7662 & T_7749;
  assign T_7751 = T_7746 | T_7748;
  assign T_7752 = T_7751 | T_7750;
  assign data_hazard_wb = wb_ctrl_wxd & T_7752;
  assign T_7754 = io_fpu_dec_ren1 & T_7745;
  assign T_7756 = io_fpu_dec_ren2 & T_7747;
  assign T_7757 = id_raddr3 == wb_waddr;
  assign T_7758 = io_fpu_dec_ren3 & T_7757;
  assign T_7760 = io_fpu_dec_wen & T_7749;
  assign T_7761 = T_7754 | T_7756;
  assign T_7762 = T_7761 | T_7758;
  assign T_7763 = T_7762 | T_7760;
  assign fp_data_hazard_wb = wb_ctrl_wfd & T_7763;
  assign T_7764 = data_hazard_wb & wb_set_sboard;
  assign T_7765 = T_7764 | fp_data_hazard_wb;
  assign id_wb_hazard = wb_reg_valid & T_7765;
  assign T_7769 = io_dmem_req_valid | dcache_blocked;
  assign T_7770 = T_7338 & T_7769;
  assign T_7773 = wb_reg_xcpt == 1'h0;
  assign T_7776 = T_7773 & T_7621;
  assign T_7777 = io_rocc_cmd_valid | rocc_blocked;
  assign T_7778 = T_7776 & T_7777;
  assign T_7779 = id_ex_hazard | id_mem_hazard;
  assign T_7780 = T_7779 | id_wb_hazard;
  assign T_7781 = T_7780 | id_sboard_hazard;
  assign T_7784 = id_ctrl_mem & dcache_blocked;
  assign T_7785 = T_7781 | T_7784;
  assign T_7786 = id_ctrl_rocc & rocc_blocked;
  assign T_7787 = T_7785 | T_7786;
  assign T_7788 = T_7787 | T_7130;
  assign ctrl_stalld = T_7788 | csr_io_csr_stall;
  assign T_7790 = io_imem_resp_valid == 1'h0;
  assign T_7791 = T_7790 | io_imem_resp_bits_replay;
  assign T_7792 = T_7791 | take_pc_mem_wb;
  assign T_7793 = T_7792 | ctrl_stalld;
  assign T_7794 = T_7793 | csr_io_interrupt;
  assign T_7797 = wb_xcpt | csr_io_eret;
  assign T_7798 = replay_wb ? wb_reg_pc : mem_npc;
  assign T_7799 = T_7797 ? csr_io_evec : T_7798;
  assign T_7800 = wb_reg_valid & wb_ctrl_fence_i;
  assign T_7802 = io_dmem_s2_nack == 1'h0;
  assign T_7803 = T_7800 & T_7802;
  assign T_7805 = ctrl_stalld == 1'h0;
  assign T_7806 = T_7805 | csr_io_interrupt;
  assign T_7807 = T_7806 | take_pc_mem;
  assign T_7810 = mem_reg_valid & T_7531;
  assign T_7811 = T_7810 & mem_wrong_npc;
  assign T_7812 = T_7811 & mem_misprediction;
  assign T_7815 = T_7812 & T_7604;
  assign T_7816 = mem_ctrl_jal | mem_ctrl_jalr;
  assign T_7817 = mem_reg_inst[19:15];
  assign T_7820 = T_7817 & 5'h19;
  assign T_7821 = 5'h1 == T_7820;
  assign T_7822 = mem_ctrl_jalr & T_7821;
  assign T_7823 = mem_reg_valid & mem_ctrl_branch;
  assign T_7826 = T_7823 & T_7604;
  assign T_7827 = mem_reg_valid & io_imem_btb_update_bits_isJump;
  assign T_7830 = T_7827 & T_7531;
  assign T_7833 = T_7830 & T_7604;
  assign T_7834 = mem_waddr[0];
  assign T_7835 = mem_ctrl_wxd & T_7834;
  assign T_7838 = T_7281 & id_ctrl_fp;
  assign T_7839 = dmem_resp_valid & T_7624;
  assign T_7840 = ex_reg_valid & ex_ctrl_mem;
  assign ex_dcache_tag = {ex_waddr,ex_ctrl_fp};
  assign T_7843 = mem_ctrl_fp ? io_fpu_store_data : {{32'd0}, mem_reg_rs2};
  assign T_7846 = replay_wb_common == 1'h0;
  assign T_7847 = T_7119 & T_7846;
  assign T_7850 = wb_xcpt & T_7107;
  assign T_7869_funct = T_7887;
  assign T_7869_rs2 = T_7886;
  assign T_7869_rs1 = T_7885;
  assign T_7869_xd = T_7884;
  assign T_7869_xs1 = T_7883;
  assign T_7869_xs2 = T_7882;
  assign T_7869_rd = T_7881;
  assign T_7869_opcode = T_7880;
  assign T_7879 = wb_reg_inst;
  assign T_7880 = T_7879[6:0];
  assign T_7881 = T_7879[11:7];
  assign T_7882 = T_7879[12];
  assign T_7883 = T_7879[13];
  assign T_7884 = T_7879[14];
  assign T_7885 = T_7879[19:15];
  assign T_7886 = T_7879[24:20];
  assign T_7887 = T_7879[31:25];
  assign T_7888 = csr_io_time;
  assign T_7890 = rf_wen ? rf_waddr : 8'h0;
  assign T_7891 = wb_reg_inst[19:15];
  assign T_7894 = wb_reg_inst[24:20];
  assign T_7898 = reset == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_271 = {1{$random}};
  ex_ctrl_legal = GEN_271[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_272 = {1{$random}};
  ex_ctrl_fp = GEN_272[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_273 = {1{$random}};
  ex_ctrl_rocc = GEN_273[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_274 = {1{$random}};
  ex_ctrl_branch = GEN_274[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_275 = {1{$random}};
  ex_ctrl_jal = GEN_275[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_276 = {1{$random}};
  ex_ctrl_jalr = GEN_276[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_277 = {1{$random}};
  ex_ctrl_rxs2 = GEN_277[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_278 = {1{$random}};
  ex_ctrl_rxs1 = GEN_278[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_279 = {1{$random}};
  ex_ctrl_sel_alu2 = GEN_279[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_280 = {1{$random}};
  ex_ctrl_sel_alu1 = GEN_280[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_281 = {1{$random}};
  ex_ctrl_sel_imm = GEN_281[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_282 = {1{$random}};
  ex_ctrl_alu_dw = GEN_282[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_283 = {1{$random}};
  ex_ctrl_alu_fn = GEN_283[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_284 = {1{$random}};
  ex_ctrl_mem = GEN_284[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_285 = {1{$random}};
  ex_ctrl_mem_cmd = GEN_285[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_286 = {1{$random}};
  ex_ctrl_mem_type = GEN_286[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_287 = {1{$random}};
  ex_ctrl_rfs1 = GEN_287[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_288 = {1{$random}};
  ex_ctrl_rfs2 = GEN_288[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_289 = {1{$random}};
  ex_ctrl_rfs3 = GEN_289[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_290 = {1{$random}};
  ex_ctrl_wfd = GEN_290[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_291 = {1{$random}};
  ex_ctrl_div = GEN_291[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_292 = {1{$random}};
  ex_ctrl_wxd = GEN_292[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_293 = {1{$random}};
  ex_ctrl_csr = GEN_293[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_294 = {1{$random}};
  ex_ctrl_fence_i = GEN_294[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_295 = {1{$random}};
  ex_ctrl_fence = GEN_295[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_296 = {1{$random}};
  ex_ctrl_amo = GEN_296[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_297 = {1{$random}};
  mem_ctrl_legal = GEN_297[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_298 = {1{$random}};
  mem_ctrl_fp = GEN_298[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_299 = {1{$random}};
  mem_ctrl_rocc = GEN_299[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_300 = {1{$random}};
  mem_ctrl_branch = GEN_300[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_301 = {1{$random}};
  mem_ctrl_jal = GEN_301[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_302 = {1{$random}};
  mem_ctrl_jalr = GEN_302[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_303 = {1{$random}};
  mem_ctrl_rxs2 = GEN_303[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_304 = {1{$random}};
  mem_ctrl_rxs1 = GEN_304[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_305 = {1{$random}};
  mem_ctrl_sel_alu2 = GEN_305[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_306 = {1{$random}};
  mem_ctrl_sel_alu1 = GEN_306[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_307 = {1{$random}};
  mem_ctrl_sel_imm = GEN_307[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_308 = {1{$random}};
  mem_ctrl_alu_dw = GEN_308[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_309 = {1{$random}};
  mem_ctrl_alu_fn = GEN_309[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_310 = {1{$random}};
  mem_ctrl_mem = GEN_310[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_311 = {1{$random}};
  mem_ctrl_mem_cmd = GEN_311[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_312 = {1{$random}};
  mem_ctrl_mem_type = GEN_312[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_313 = {1{$random}};
  mem_ctrl_rfs1 = GEN_313[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_314 = {1{$random}};
  mem_ctrl_rfs2 = GEN_314[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_315 = {1{$random}};
  mem_ctrl_rfs3 = GEN_315[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_316 = {1{$random}};
  mem_ctrl_wfd = GEN_316[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_317 = {1{$random}};
  mem_ctrl_div = GEN_317[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_318 = {1{$random}};
  mem_ctrl_wxd = GEN_318[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_319 = {1{$random}};
  mem_ctrl_csr = GEN_319[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_320 = {1{$random}};
  mem_ctrl_fence_i = GEN_320[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_321 = {1{$random}};
  mem_ctrl_fence = GEN_321[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_322 = {1{$random}};
  mem_ctrl_amo = GEN_322[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_323 = {1{$random}};
  wb_ctrl_legal = GEN_323[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_324 = {1{$random}};
  wb_ctrl_fp = GEN_324[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_325 = {1{$random}};
  wb_ctrl_rocc = GEN_325[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_326 = {1{$random}};
  wb_ctrl_branch = GEN_326[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_327 = {1{$random}};
  wb_ctrl_jal = GEN_327[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_328 = {1{$random}};
  wb_ctrl_jalr = GEN_328[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_329 = {1{$random}};
  wb_ctrl_rxs2 = GEN_329[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_330 = {1{$random}};
  wb_ctrl_rxs1 = GEN_330[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_331 = {1{$random}};
  wb_ctrl_sel_alu2 = GEN_331[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_332 = {1{$random}};
  wb_ctrl_sel_alu1 = GEN_332[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_333 = {1{$random}};
  wb_ctrl_sel_imm = GEN_333[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_334 = {1{$random}};
  wb_ctrl_alu_dw = GEN_334[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_335 = {1{$random}};
  wb_ctrl_alu_fn = GEN_335[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_336 = {1{$random}};
  wb_ctrl_mem = GEN_336[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_337 = {1{$random}};
  wb_ctrl_mem_cmd = GEN_337[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_338 = {1{$random}};
  wb_ctrl_mem_type = GEN_338[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_339 = {1{$random}};
  wb_ctrl_rfs1 = GEN_339[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_340 = {1{$random}};
  wb_ctrl_rfs2 = GEN_340[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_341 = {1{$random}};
  wb_ctrl_rfs3 = GEN_341[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_342 = {1{$random}};
  wb_ctrl_wfd = GEN_342[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_343 = {1{$random}};
  wb_ctrl_div = GEN_343[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_344 = {1{$random}};
  wb_ctrl_wxd = GEN_344[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_345 = {1{$random}};
  wb_ctrl_csr = GEN_345[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_346 = {1{$random}};
  wb_ctrl_fence_i = GEN_346[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_347 = {1{$random}};
  wb_ctrl_fence = GEN_347[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_348 = {1{$random}};
  wb_ctrl_amo = GEN_348[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_349 = {1{$random}};
  ex_reg_xcpt_interrupt = GEN_349[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_350 = {1{$random}};
  ex_reg_valid = GEN_350[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_351 = {1{$random}};
  ex_reg_btb_hit = GEN_351[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_352 = {1{$random}};
  ex_reg_btb_resp_taken = GEN_352[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_353 = {1{$random}};
  ex_reg_btb_resp_mask = GEN_353[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_354 = {1{$random}};
  ex_reg_btb_resp_bridx = GEN_354[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_355 = {1{$random}};
  ex_reg_btb_resp_target = GEN_355[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_356 = {1{$random}};
  ex_reg_btb_resp_entry = GEN_356[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_357 = {1{$random}};
  ex_reg_btb_resp_bht_history = GEN_357[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_358 = {1{$random}};
  ex_reg_btb_resp_bht_value = GEN_358[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_359 = {1{$random}};
  ex_reg_xcpt = GEN_359[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_360 = {1{$random}};
  ex_reg_flush_pipe = GEN_360[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_361 = {1{$random}};
  ex_reg_load_use = GEN_361[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_362 = {1{$random}};
  ex_reg_cause = GEN_362[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_363 = {1{$random}};
  ex_reg_replay = GEN_363[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_364 = {1{$random}};
  ex_reg_pc = GEN_364[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_365 = {1{$random}};
  ex_reg_inst = GEN_365[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_366 = {1{$random}};
  mem_reg_xcpt_interrupt = GEN_366[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_367 = {1{$random}};
  mem_reg_valid = GEN_367[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_368 = {1{$random}};
  mem_reg_btb_hit = GEN_368[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_369 = {1{$random}};
  mem_reg_btb_resp_taken = GEN_369[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_370 = {1{$random}};
  mem_reg_btb_resp_mask = GEN_370[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_371 = {1{$random}};
  mem_reg_btb_resp_bridx = GEN_371[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_372 = {1{$random}};
  mem_reg_btb_resp_target = GEN_372[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_373 = {1{$random}};
  mem_reg_btb_resp_entry = GEN_373[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_374 = {1{$random}};
  mem_reg_btb_resp_bht_history = GEN_374[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_375 = {1{$random}};
  mem_reg_btb_resp_bht_value = GEN_375[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_376 = {1{$random}};
  mem_reg_xcpt = GEN_376[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_377 = {1{$random}};
  mem_reg_replay = GEN_377[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_378 = {1{$random}};
  mem_reg_flush_pipe = GEN_378[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_379 = {1{$random}};
  mem_reg_cause = GEN_379[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_380 = {1{$random}};
  mem_reg_slow_bypass = GEN_380[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_381 = {1{$random}};
  mem_reg_load = GEN_381[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_382 = {1{$random}};
  mem_reg_store = GEN_382[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_383 = {1{$random}};
  mem_reg_pc = GEN_383[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_384 = {1{$random}};
  mem_reg_inst = GEN_384[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_385 = {1{$random}};
  mem_reg_wdata = GEN_385[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_386 = {1{$random}};
  mem_reg_rs2 = GEN_386[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_387 = {1{$random}};
  wb_reg_valid = GEN_387[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_388 = {1{$random}};
  wb_reg_xcpt = GEN_388[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_389 = {1{$random}};
  wb_reg_mem_xcpt = GEN_389[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_390 = {1{$random}};
  wb_reg_replay = GEN_390[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_391 = {1{$random}};
  wb_reg_cause = GEN_391[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_392 = {1{$random}};
  wb_reg_pc = GEN_392[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_393 = {1{$random}};
  wb_reg_inst = GEN_393[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_394 = {1{$random}};
  wb_reg_wdata = GEN_394[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_395 = {1{$random}};
  wb_reg_rs2 = GEN_395[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_396 = {1{$random}};
  id_reg_fence = GEN_396[0:0];
  `endif
  GEN_397 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 31; initvar = initvar+1)
    T_6999[initvar] = GEN_397[31:0];
  `endif
  GEN_398 = {1{$random}};
  GEN_399 = {1{$random}};
  `ifdef RANDOMIZE
  GEN_400 = {1{$random}};
  ex_reg_rs_bypass_0 = GEN_400[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_401 = {1{$random}};
  ex_reg_rs_bypass_1 = GEN_401[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_402 = {1{$random}};
  ex_reg_rs_lsb_0 = GEN_402[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_403 = {1{$random}};
  ex_reg_rs_lsb_1 = GEN_403[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_404 = {1{$random}};
  ex_reg_rs_msb_0 = GEN_404[29:0];
  `endif
  `ifdef RANDOMIZE
  GEN_405 = {1{$random}};
  ex_reg_rs_msb_1 = GEN_405[29:0];
  `endif
  `ifdef RANDOMIZE
  GEN_406 = {1{$random}};
  T_7598 = GEN_406[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_407 = {1{$random}};
  T_7664 = GEN_407[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_408 = {1{$random}};
  dcache_blocked = GEN_408[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_409 = {1{$random}};
  rocc_blocked = GEN_409[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_410 = {1{$random}};
  T_7892 = GEN_410[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_411 = {1{$random}};
  T_7893 = GEN_411[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_412 = {1{$random}};
  T_7895 = GEN_412[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_413 = {1{$random}};
  T_7896 = GEN_413[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_414 = {1{$random}};
  GEN_154 = GEN_414[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_415 = {1{$random}};
  GEN_155 = GEN_415[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_416 = {1{$random}};
  GEN_156 = GEN_416[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_417 = {1{$random}};
  GEN_157 = GEN_417[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_418 = {1{$random}};
  GEN_158 = GEN_418[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_419 = {1{$random}};
  GEN_161 = GEN_419[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_420 = {1{$random}};
  GEN_162 = GEN_420[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_421 = {1{$random}};
  GEN_164 = GEN_421[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_422 = {1{$random}};
  GEN_165 = GEN_422[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_423 = {1{$random}};
  GEN_174 = GEN_423[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_424 = {1{$random}};
  GEN_175 = GEN_424[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_425 = {1{$random}};
  GEN_176 = GEN_425[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_426 = {1{$random}};
  GEN_177 = GEN_426[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_427 = {1{$random}};
  GEN_178 = GEN_427[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_428 = {1{$random}};
  GEN_179 = GEN_428[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_429 = {1{$random}};
  GEN_180 = GEN_429[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_430 = {1{$random}};
  GEN_181 = GEN_430[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_431 = {1{$random}};
  GEN_182 = GEN_431[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_432 = {1{$random}};
  GEN_183 = GEN_432[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_433 = {1{$random}};
  GEN_184 = GEN_433[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_434 = {1{$random}};
  GEN_185 = GEN_434[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_435 = {1{$random}};
  GEN_186 = GEN_435[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_436 = {3{$random}};
  GEN_187 = GEN_436[64:0];
  `endif
  `ifdef RANDOMIZE
  GEN_437 = {3{$random}};
  GEN_188 = GEN_437[64:0];
  `endif
  `ifdef RANDOMIZE
  GEN_438 = {3{$random}};
  GEN_189 = GEN_438[64:0];
  `endif
  `ifdef RANDOMIZE
  GEN_439 = {1{$random}};
  GEN_190 = GEN_439[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_440 = {1{$random}};
  GEN_191 = GEN_440[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_441 = {1{$random}};
  GEN_192 = GEN_441[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_442 = {1{$random}};
  GEN_193 = GEN_442[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_443 = {1{$random}};
  GEN_194 = GEN_443[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_444 = {1{$random}};
  GEN_195 = GEN_444[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_445 = {1{$random}};
  GEN_196 = GEN_445[8:0];
  `endif
  `ifdef RANDOMIZE
  GEN_446 = {1{$random}};
  GEN_197 = GEN_446[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_447 = {1{$random}};
  GEN_198 = GEN_447[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_448 = {1{$random}};
  GEN_199 = GEN_448[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_449 = {1{$random}};
  GEN_200 = GEN_449[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_450 = {1{$random}};
  GEN_201 = GEN_450[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_451 = {1{$random}};
  GEN_202 = GEN_451[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_452 = {1{$random}};
  GEN_203 = GEN_452[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_453 = {1{$random}};
  GEN_204 = GEN_453[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_454 = {1{$random}};
  GEN_205 = GEN_454[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_455 = {1{$random}};
  GEN_206 = GEN_455[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_456 = {1{$random}};
  GEN_207 = GEN_456[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_457 = {1{$random}};
  GEN_208 = GEN_457[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_458 = {1{$random}};
  GEN_209 = GEN_458[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_459 = {1{$random}};
  GEN_210 = GEN_459[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_460 = {1{$random}};
  GEN_211 = GEN_460[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_461 = {1{$random}};
  GEN_212 = GEN_461[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_462 = {1{$random}};
  GEN_213 = GEN_462[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_463 = {1{$random}};
  GEN_214 = GEN_463[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_464 = {1{$random}};
  GEN_215 = GEN_464[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_465 = {1{$random}};
  GEN_216 = GEN_465[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_466 = {2{$random}};
  GEN_217 = GEN_466[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_467 = {1{$random}};
  GEN_218 = GEN_467[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_468 = {1{$random}};
  GEN_219 = GEN_468[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_469 = {3{$random}};
  GEN_220 = GEN_469[64:0];
  `endif
  `ifdef RANDOMIZE
  GEN_470 = {1{$random}};
  GEN_221 = GEN_470[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_471 = {1{$random}};
  GEN_222 = GEN_471[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_472 = {1{$random}};
  GEN_223 = GEN_472[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_473 = {1{$random}};
  GEN_224 = GEN_473[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_474 = {1{$random}};
  GEN_225 = GEN_474[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_475 = {1{$random}};
  GEN_226 = GEN_475[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_476 = {1{$random}};
  GEN_227 = GEN_476[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_477 = {1{$random}};
  GEN_228 = GEN_477[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_478 = {1{$random}};
  GEN_229 = GEN_478[8:0];
  `endif
  `ifdef RANDOMIZE
  GEN_479 = {1{$random}};
  GEN_230 = GEN_479[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_480 = {1{$random}};
  GEN_231 = GEN_480[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_481 = {1{$random}};
  GEN_232 = GEN_481[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_482 = {1{$random}};
  GEN_233 = GEN_482[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_483 = {1{$random}};
  GEN_234 = GEN_483[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_484 = {1{$random}};
  GEN_235 = GEN_484[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_485 = {1{$random}};
  GEN_236 = GEN_485[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_486 = {1{$random}};
  GEN_237 = GEN_486[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_487 = {1{$random}};
  GEN_238 = GEN_487[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_488 = {1{$random}};
  GEN_239 = GEN_488[25:0];
  `endif
  `ifdef RANDOMIZE
  GEN_489 = {1{$random}};
  GEN_240 = GEN_489[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_490 = {1{$random}};
  GEN_241 = GEN_490[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_491 = {1{$random}};
  GEN_242 = GEN_491[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_492 = {1{$random}};
  GEN_243 = GEN_492[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_493 = {1{$random}};
  GEN_244 = GEN_493[11:0];
  `endif
  `ifdef RANDOMIZE
  GEN_494 = {2{$random}};
  GEN_245 = GEN_494[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_495 = {1{$random}};
  GEN_246 = GEN_495[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_496 = {1{$random}};
  GEN_247 = GEN_496[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_497 = {1{$random}};
  GEN_248 = GEN_497[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_498 = {1{$random}};
  GEN_249 = GEN_498[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_499 = {1{$random}};
  GEN_250 = GEN_499[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_500 = {1{$random}};
  GEN_251 = GEN_500[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_501 = {1{$random}};
  GEN_252 = GEN_501[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_502 = {1{$random}};
  GEN_253 = GEN_502[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_503 = {1{$random}};
  GEN_254 = GEN_503[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_504 = {1{$random}};
  GEN_255 = GEN_504[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_505 = {1{$random}};
  GEN_256 = GEN_505[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_506 = {1{$random}};
  GEN_257 = GEN_506[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_507 = {1{$random}};
  GEN_258 = GEN_507[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_508 = {1{$random}};
  GEN_259 = GEN_508[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_509 = {1{$random}};
  GEN_260 = GEN_509[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_510 = {1{$random}};
  GEN_261 = GEN_510[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_511 = {1{$random}};
  GEN_262 = GEN_511[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_512 = {1{$random}};
  GEN_263 = GEN_512[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_513 = {1{$random}};
  GEN_264 = GEN_513[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_514 = {1{$random}};
  GEN_265 = GEN_514[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_515 = {1{$random}};
  GEN_266 = GEN_515[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_516 = {3{$random}};
  GEN_267 = GEN_516[64:0];
  `endif
  `ifdef RANDOMIZE
  GEN_517 = {3{$random}};
  GEN_268 = GEN_517[64:0];
  `endif
  `ifdef RANDOMIZE
  GEN_518 = {3{$random}};
  GEN_269 = GEN_518[64:0];
  `endif
  `ifdef RANDOMIZE
  GEN_519 = {1{$random}};
  GEN_270 = GEN_519[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_legal <= id_ctrl_legal;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_fp <= id_ctrl_fp;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_rocc <= id_ctrl_rocc;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_branch <= id_ctrl_branch;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_jal <= id_ctrl_jal;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_jalr <= id_ctrl_jalr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_rxs2 <= id_ctrl_rxs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_rxs1 <= id_ctrl_rxs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_sel_alu2 <= id_ctrl_sel_alu2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_sel_alu1 <= id_ctrl_sel_alu1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_sel_imm <= id_ctrl_sel_imm;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_alu_dw <= id_ctrl_alu_dw;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_alu_fn <= id_ctrl_alu_fn;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_mem <= id_ctrl_mem;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_mem_cmd <= id_ctrl_mem_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_mem_type <= id_ctrl_mem_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_rfs1 <= id_ctrl_rfs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_rfs2 <= id_ctrl_rfs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_rfs3 <= id_ctrl_rfs3;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_wfd <= id_ctrl_wfd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_div <= id_ctrl_div;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_wxd <= id_ctrl_wxd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        if(id_csr_ren) begin
          ex_ctrl_csr <= 3'h5;
        end else begin
          ex_ctrl_csr <= id_ctrl_csr;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        if(T_7297) begin
          ex_ctrl_fence_i <= 1'h1;
        end else begin
          ex_ctrl_fence_i <= id_ctrl_fence_i;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_fence <= id_ctrl_fence;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_ctrl_amo <= id_ctrl_amo;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_legal <= ex_ctrl_legal;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_fp <= ex_ctrl_fp;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rocc <= ex_ctrl_rocc;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_branch <= ex_ctrl_branch;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_jal <= ex_ctrl_jal;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_jalr <= ex_ctrl_jalr;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rxs2 <= ex_ctrl_rxs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rxs1 <= ex_ctrl_rxs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_sel_alu2 <= ex_ctrl_sel_alu2;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_sel_alu1 <= ex_ctrl_sel_alu1;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_sel_imm <= ex_ctrl_sel_imm;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_alu_dw <= ex_ctrl_alu_dw;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_alu_fn <= ex_ctrl_alu_fn;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_mem <= ex_ctrl_mem;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_mem_cmd <= ex_ctrl_mem_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_mem_type <= ex_ctrl_mem_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rfs1 <= ex_ctrl_rfs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rfs2 <= ex_ctrl_rfs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_rfs3 <= ex_ctrl_rfs3;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_wfd <= ex_ctrl_wfd;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_div <= ex_ctrl_div;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_wxd <= ex_ctrl_wxd;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_csr <= ex_ctrl_csr;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_fence_i <= ex_ctrl_fence_i;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_fence <= ex_ctrl_fence;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_ctrl_amo <= ex_ctrl_amo;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_legal <= mem_ctrl_legal;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_fp <= mem_ctrl_fp;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_rocc <= mem_ctrl_rocc;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_branch <= mem_ctrl_branch;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_jal <= mem_ctrl_jal;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_jalr <= mem_ctrl_jalr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_rxs2 <= mem_ctrl_rxs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_rxs1 <= mem_ctrl_rxs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_sel_alu2 <= mem_ctrl_sel_alu2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_sel_alu1 <= mem_ctrl_sel_alu1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_sel_imm <= mem_ctrl_sel_imm;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_alu_dw <= mem_ctrl_alu_dw;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_alu_fn <= mem_ctrl_alu_fn;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_mem <= mem_ctrl_mem;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_mem_cmd <= mem_ctrl_mem_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_mem_type <= mem_ctrl_mem_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_rfs1 <= mem_ctrl_rfs1;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_rfs2 <= mem_ctrl_rfs2;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_rfs3 <= mem_ctrl_rfs3;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_wfd <= mem_ctrl_wfd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_div <= mem_ctrl_div;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_wxd <= mem_ctrl_wxd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_csr <= mem_ctrl_csr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_fence_i <= mem_ctrl_fence_i;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_fence <= mem_ctrl_fence;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_ctrl_amo <= mem_ctrl_amo;
      end
    end
    if(1'h0) begin
    end else begin
      ex_reg_xcpt_interrupt <= T_7292;
    end
    if(1'h0) begin
    end else begin
      ex_reg_valid <= T_7281;
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_reg_btb_hit <= io_imem_btb_resp_valid;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        if(io_imem_btb_resp_valid) begin
          ex_reg_btb_resp_taken <= io_imem_btb_resp_bits_taken;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        if(io_imem_btb_resp_valid) begin
          ex_reg_btb_resp_mask <= io_imem_btb_resp_bits_mask;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        if(io_imem_btb_resp_valid) begin
          ex_reg_btb_resp_bridx <= io_imem_btb_resp_bits_bridx;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        if(io_imem_btb_resp_valid) begin
          ex_reg_btb_resp_target <= io_imem_btb_resp_bits_target;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        if(io_imem_btb_resp_valid) begin
          ex_reg_btb_resp_entry <= io_imem_btb_resp_bits_entry;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        if(io_imem_btb_resp_valid) begin
          ex_reg_btb_resp_bht_history <= io_imem_btb_resp_bits_bht_history;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        if(io_imem_btb_resp_valid) begin
          ex_reg_btb_resp_bht_value <= io_imem_btb_resp_bits_bht_value;
        end
      end
    end
    if(1'h0) begin
    end else begin
      ex_reg_xcpt <= T_7288;
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        if(T_7297) begin
          ex_reg_flush_pipe <= 1'h1;
        end else begin
          ex_reg_flush_pipe <= T_7296;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_reg_load_use <= id_load_use;
      end
    end
    if(1'h0) begin
    end else begin
      if(id_xcpt) begin
        if(csr_io_interrupt) begin
          ex_reg_cause <= csr_io_interrupt_cause;
        end else begin
          ex_reg_cause <= {{30'd0}, T_7137};
        end
      end
    end
    if(1'h0) begin
    end else begin
      ex_reg_replay <= T_7285;
    end
    if(1'h0) begin
    end else begin
      if(T_7333) begin
        ex_reg_pc <= io_imem_resp_bits_pc;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7333) begin
        ex_reg_inst <= io_imem_resp_bits_data_0;
      end
    end
    if(1'h0) begin
    end else begin
      mem_reg_xcpt_interrupt <= T_7543;
    end
    if(1'h0) begin
    end else begin
      mem_reg_valid <= T_7534;
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_btb_hit <= ex_reg_btb_hit;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_taken <= ex_reg_btb_resp_taken;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_mask <= ex_reg_btb_resp_mask;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_bridx <= ex_reg_btb_resp_bridx;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_target <= ex_reg_btb_resp_target;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_entry <= ex_reg_btb_resp_entry;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_bht_history <= ex_reg_btb_resp_bht_history;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(ex_reg_btb_hit) begin
          mem_reg_btb_resp_bht_value <= ex_reg_btb_resp_bht_value;
        end
      end
    end
    if(1'h0) begin
    end else begin
      mem_reg_xcpt <= T_7540;
    end
    if(1'h0) begin
    end else begin
      mem_reg_replay <= T_7537;
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_flush_pipe <= ex_reg_flush_pipe;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_xcpt) begin
        if(T_7365) begin
          mem_reg_cause <= ex_reg_cause;
        end else begin
          mem_reg_cause <= 32'h2;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_slow_bypass <= ex_slow_bypass;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_load <= T_7553;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_store <= T_7561;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_pc <= ex_reg_pc;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_inst <= ex_reg_inst;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        mem_reg_wdata <= alu_io_out;
      end
    end
    if(1'h0) begin
    end else begin
      if(ex_pc_valid) begin
        if(T_7563) begin
          if(ex_reg_rs_bypass_1) begin
            mem_reg_rs2 <= GEN_1;
          end else begin
            mem_reg_rs2 <= T_7192;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      wb_reg_valid <= T_7602;
    end
    if(1'h0) begin
    end else begin
      wb_reg_xcpt <= T_7608;
    end
    if(1'h0) begin
    end else begin
      wb_reg_mem_xcpt <= T_7613;
    end
    if(1'h0) begin
    end else begin
      wb_reg_replay <= T_7605;
    end
    if(1'h0) begin
    end else begin
      if(mem_xcpt) begin
        if(T_7588) begin
          wb_reg_cause <= mem_reg_cause;
        end else begin
          wb_reg_cause <= {{29'd0}, mem_new_cause};
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_reg_pc <= mem_reg_pc;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        wb_reg_inst <= mem_reg_inst;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        if(T_7616) begin
          wb_reg_wdata <= io_fpu_toint_data;
        end else begin
          wb_reg_wdata <= mem_int_wdata;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7615) begin
        if(mem_ctrl_rocc) begin
          wb_reg_rs2 <= mem_reg_rs2;
        end
      end
    end
    if(reset) begin
      id_reg_fence <= 1'h0;
    end else begin
      id_reg_fence <= T_7122;
    end
    if(T_6999_T_7648_en & T_6999_T_7648_mask) begin
      T_6999[T_6999_T_7648_addr] <= T_6999_T_7648_data;
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_reg_rs_bypass_0 <= T_7302;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        ex_reg_rs_bypass_1 <= T_7317;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        if(T_7312) begin
          ex_reg_rs_lsb_0 <= T_7313;
        end else begin
          if(T_7147) begin
            ex_reg_rs_lsb_0 <= 2'h0;
          end else begin
            if(T_7150) begin
              ex_reg_rs_lsb_0 <= 2'h1;
            end else begin
              if(T_7152) begin
                ex_reg_rs_lsb_0 <= 2'h2;
              end else begin
                ex_reg_rs_lsb_0 <= 2'h3;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        if(T_7327) begin
          ex_reg_rs_lsb_1 <= T_7328;
        end else begin
          if(T_7155) begin
            ex_reg_rs_lsb_1 <= 2'h0;
          end else begin
            if(T_7158) begin
              ex_reg_rs_lsb_1 <= 2'h1;
            end else begin
              if(T_7160) begin
                ex_reg_rs_lsb_1 <= 2'h2;
              end else begin
                ex_reg_rs_lsb_1 <= 2'h3;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        if(T_7312) begin
          ex_reg_rs_msb_0 <= T_7314;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_7281) begin
        if(T_7327) begin
          ex_reg_rs_msb_1 <= T_7329;
        end
      end
    end
    if(1'h0) begin
    end else begin
      T_7598 <= T_7597;
    end
    if(reset) begin
      T_7664 <= 32'h0;
    end else begin
      T_7664 <= GEN_169[31:0];
    end
    if(1'h0) begin
    end else begin
      dcache_blocked <= T_7770;
    end
    if(1'h0) begin
    end else begin
      rocc_blocked <= T_7778;
    end
    if(1'h0) begin
    end else begin
      if(ex_reg_rs_bypass_0) begin
        T_7892 <= GEN_0;
      end else begin
        T_7892 <= T_7190;
      end
    end
    if(1'h0) begin
    end else begin
      T_7893 <= T_7892;
    end
    if(1'h0) begin
    end else begin
      if(ex_reg_rs_bypass_1) begin
        T_7895 <= GEN_1;
      end else begin
        T_7895 <= T_7192;
      end
    end
    if(1'h0) begin
    end else begin
      T_7896 <= T_7895;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_7898) begin
          $fwrite(32'h80000002,"C%d: %d [%d] pc=[%h] W[r%d=%h][%d] R[r%d=%h] R[r%d=%h] inst=[%h] DASM(%h)\n",io_prci_id,T_7888,wb_valid,wb_reg_pc,T_7890,rf_wdata,rf_wen,T_7891,T_7893,T_7894,T_7896,wb_reg_inst,wb_reg_inst);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module FlowThroughSerializer(
  input   clk,
  input   reset,
  output  io_in_ready,
  input   io_in_valid,
  input  [2:0] io_in_bits_addr_beat,
  input   io_in_bits_client_xact_id,
  input  [1:0] io_in_bits_manager_xact_id,
  input   io_in_bits_is_builtin_type,
  input  [3:0] io_in_bits_g_type,
  input  [63:0] io_in_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output  io_out_bits_client_xact_id,
  output [1:0] io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_cnt,
  output  io_done
);
  assign io_in_ready = io_out_ready;
  assign io_out_valid = io_in_valid;
  assign io_out_bits_addr_beat = io_in_bits_addr_beat;
  assign io_out_bits_client_xact_id = io_in_bits_client_xact_id;
  assign io_out_bits_manager_xact_id = io_in_bits_manager_xact_id;
  assign io_out_bits_is_builtin_type = io_in_bits_is_builtin_type;
  assign io_out_bits_g_type = io_in_bits_g_type;
  assign io_out_bits_data = io_in_bits_data;
  assign io_cnt = 1'h0;
  assign io_done = 1'h1;
endmodule
module ICache(
  input   clk,
  input   reset,
  input   io_req_valid,
  input  [31:0] io_req_bits_addr,
  input  [19:0] io_s1_ppn,
  input   io_s1_kill,
  input   io_s2_kill,
  input   io_resp_ready,
  output  io_resp_valid,
  output [31:0] io_resp_bits_data,
  output [63:0] io_resp_bits_datablock,
  input   io_invalidate,
  input   io_mem_acquire_ready,
  output  io_mem_acquire_valid,
  output [25:0] io_mem_acquire_bits_addr_block,
  output  io_mem_acquire_bits_client_xact_id,
  output [2:0] io_mem_acquire_bits_addr_beat,
  output  io_mem_acquire_bits_is_builtin_type,
  output [2:0] io_mem_acquire_bits_a_type,
  output [11:0] io_mem_acquire_bits_union,
  output [63:0] io_mem_acquire_bits_data,
  output  io_mem_grant_ready,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input   io_mem_grant_bits_client_xact_id,
  input  [1:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data
);
  reg [1:0] state;
  reg [31:0] GEN_4;
  reg  invalidated;
  reg [31:0] GEN_5;
  wire  stall;
  wire  rdy;
  reg [31:0] refill_addr;
  reg [31:0] GEN_6;
  wire  s1_any_tag_hit;
  reg  s1_valid;
  reg [31:0] GEN_7;
  reg [31:0] s1_vaddr;
  reg [31:0] GEN_8;
  wire [11:0] T_827;
  wire [31:0] s1_paddr;
  wire [18:0] s1_tag;
  wire  T_828;
  wire [31:0] s0_vaddr;
  wire  T_830;
  wire  T_833;
  wire  T_834;
  wire  T_835;
  wire [31:0] GEN_0;
  wire  T_839;
  wire  T_840;
  wire  out_valid;
  wire [6:0] s1_idx;
  wire  s1_hit;
  wire  T_842;
  wire  s1_miss;
  wire  T_845;
  wire  T_846;
  wire  T_848;
  wire [31:0] GEN_1;
  wire [18:0] refill_tag;
  wire  FlowThroughSerializer_1_clk;
  wire  FlowThroughSerializer_1_reset;
  wire  FlowThroughSerializer_1_io_in_ready;
  wire  FlowThroughSerializer_1_io_in_valid;
  wire [2:0] FlowThroughSerializer_1_io_in_bits_addr_beat;
  wire  FlowThroughSerializer_1_io_in_bits_client_xact_id;
  wire [1:0] FlowThroughSerializer_1_io_in_bits_manager_xact_id;
  wire  FlowThroughSerializer_1_io_in_bits_is_builtin_type;
  wire [3:0] FlowThroughSerializer_1_io_in_bits_g_type;
  wire [63:0] FlowThroughSerializer_1_io_in_bits_data;
  wire  FlowThroughSerializer_1_io_out_ready;
  wire  FlowThroughSerializer_1_io_out_valid;
  wire [2:0] FlowThroughSerializer_1_io_out_bits_addr_beat;
  wire  FlowThroughSerializer_1_io_out_bits_client_xact_id;
  wire [1:0] FlowThroughSerializer_1_io_out_bits_manager_xact_id;
  wire  FlowThroughSerializer_1_io_out_bits_is_builtin_type;
  wire [3:0] FlowThroughSerializer_1_io_out_bits_g_type;
  wire [63:0] FlowThroughSerializer_1_io_out_bits_data;
  wire  FlowThroughSerializer_1_io_cnt;
  wire  FlowThroughSerializer_1_io_done;
  wire  T_849;
  reg [2:0] refill_cnt;
  reg [31:0] GEN_9;
  wire  T_852;
  wire [3:0] T_854;
  wire [2:0] T_855;
  wire [2:0] GEN_2;
  wire  refill_wrap;
  wire  T_856;
  wire  refill_done;
  reg [18:0] tag_array_0 [0:127];
  reg [31:0] GEN_10;
  wire [18:0] tag_array_0_tag_rdata_data;
  wire [6:0] tag_array_0_tag_rdata_addr;
  wire  tag_array_0_tag_rdata_en;
  reg [6:0] GEN_11;
  reg [31:0] GEN_17;
  reg  GEN_18;
  reg [31:0] GEN_19;
  wire [18:0] tag_array_0_T_893_data;
  wire [6:0] tag_array_0_T_893_addr;
  wire  tag_array_0_T_893_mask;
  wire  tag_array_0_T_893_en;
  wire [6:0] T_866;
  wire [6:0] T_871;
  wire [18:0] T_880_0;
  wire  T_889_0;
  wire  GEN_12;
  reg [127:0] vb_array;
  reg [127:0] GEN_21;
  wire  T_897;
  wire  T_898;
  wire [7:0] T_899;
  wire [255:0] T_902;
  wire [255:0] GEN_36;
  wire [255:0] T_903;
  wire [127:0] T_904;
  wire [255:0] GEN_37;
  wire [255:0] T_905;
  wire [255:0] T_906;
  wire [255:0] GEN_13;
  wire [255:0] GEN_14;
  wire  GEN_15;
  wire  s1_disparity_0;
  wire  T_917;
  wire [255:0] GEN_16;
  wire  s1_tag_match_0;
  wire  s1_tag_hit_0;
  wire [63:0] s1_dout_0;
  wire  T_950;
  wire [127:0] T_954;
  wire  T_955;
  wire  T_957;
  wire [18:0] T_961;
  wire  T_962;
  wire  T_963;
  wire  T_970;
  wire  T_971;
  reg [63:0] T_974 [0:1023];
  reg [63:0] GEN_22;
  wire [63:0] T_974_T_987_data;
  wire [9:0] T_974_T_987_addr;
  wire  T_974_T_987_en;
  reg [9:0] GEN_38;
  reg [31:0] GEN_39;
  reg  GEN_42;
  reg [31:0] GEN_43;
  wire [63:0] T_974_T_980_data;
  wire [9:0] T_974_T_980_addr;
  wire  T_974_T_980_mask;
  wire  T_974_T_980_en;
  wire  T_977;
  wire [9:0] GEN_40;
  wire [9:0] T_978;
  wire [9:0] GEN_41;
  wire [9:0] T_979;
  wire [63:0] GEN_20;
  wire [9:0] T_981;
  wire [9:0] T_986;
  wire  T_989;
  reg  T_990;
  reg [31:0] GEN_44;
  wire  GEN_23;
  reg  T_995_0;
  reg [31:0] GEN_45;
  wire  GEN_24;
  reg [63:0] T_1001_0;
  reg [63:0] GEN_46;
  wire [63:0] GEN_25;
  wire  T_1003;
  wire  T_1005;
  wire  T_1006;
  wire [25:0] T_1007;
  wire [25:0] T_1110_addr_block;
  wire  T_1110_client_xact_id;
  wire [2:0] T_1110_addr_beat;
  wire  T_1110_is_builtin_type;
  wire [2:0] T_1110_a_type;
  wire [11:0] T_1110_union;
  wire [63:0] T_1110_data;
  wire  T_1138;
  wire [1:0] GEN_26;
  wire [1:0] GEN_27;
  wire  GEN_28;
  wire  T_1140;
  wire [1:0] GEN_29;
  wire [1:0] GEN_30;
  wire [1:0] GEN_31;
  wire  T_1141;
  wire [1:0] GEN_32;
  wire [1:0] GEN_33;
  wire  T_1142;
  wire [1:0] GEN_34;
  wire [1:0] GEN_35;
  reg [31:0] GEN_3;
  reg [31:0] GEN_47;
  FlowThroughSerializer FlowThroughSerializer_1 (
    .clk(FlowThroughSerializer_1_clk),
    .reset(FlowThroughSerializer_1_reset),
    .io_in_ready(FlowThroughSerializer_1_io_in_ready),
    .io_in_valid(FlowThroughSerializer_1_io_in_valid),
    .io_in_bits_addr_beat(FlowThroughSerializer_1_io_in_bits_addr_beat),
    .io_in_bits_client_xact_id(FlowThroughSerializer_1_io_in_bits_client_xact_id),
    .io_in_bits_manager_xact_id(FlowThroughSerializer_1_io_in_bits_manager_xact_id),
    .io_in_bits_is_builtin_type(FlowThroughSerializer_1_io_in_bits_is_builtin_type),
    .io_in_bits_g_type(FlowThroughSerializer_1_io_in_bits_g_type),
    .io_in_bits_data(FlowThroughSerializer_1_io_in_bits_data),
    .io_out_ready(FlowThroughSerializer_1_io_out_ready),
    .io_out_valid(FlowThroughSerializer_1_io_out_valid),
    .io_out_bits_addr_beat(FlowThroughSerializer_1_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(FlowThroughSerializer_1_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(FlowThroughSerializer_1_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(FlowThroughSerializer_1_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(FlowThroughSerializer_1_io_out_bits_g_type),
    .io_out_bits_data(FlowThroughSerializer_1_io_out_bits_data),
    .io_cnt(FlowThroughSerializer_1_io_cnt),
    .io_done(FlowThroughSerializer_1_io_done)
  );
  assign io_resp_valid = T_990;
  assign io_resp_bits_data = GEN_3;
  assign io_resp_bits_datablock = T_1001_0;
  assign io_mem_acquire_valid = T_1006;
  assign io_mem_acquire_bits_addr_block = T_1110_addr_block;
  assign io_mem_acquire_bits_client_xact_id = T_1110_client_xact_id;
  assign io_mem_acquire_bits_addr_beat = T_1110_addr_beat;
  assign io_mem_acquire_bits_is_builtin_type = T_1110_is_builtin_type;
  assign io_mem_acquire_bits_a_type = T_1110_a_type;
  assign io_mem_acquire_bits_union = T_1110_union;
  assign io_mem_acquire_bits_data = T_1110_data;
  assign io_mem_grant_ready = FlowThroughSerializer_1_io_in_ready;
  assign stall = io_resp_ready == 1'h0;
  assign rdy = T_846;
  assign s1_any_tag_hit = T_971;
  assign T_827 = s1_vaddr[11:0];
  assign s1_paddr = {io_s1_ppn,T_827};
  assign s1_tag = s1_paddr[31:13];
  assign T_828 = s1_valid & stall;
  assign s0_vaddr = T_828 ? s1_vaddr : io_req_bits_addr;
  assign T_830 = io_req_valid & rdy;
  assign T_833 = io_s1_kill == 1'h0;
  assign T_834 = T_828 & T_833;
  assign T_835 = T_830 | T_834;
  assign GEN_0 = T_830 ? io_req_bits_addr : s1_vaddr;
  assign T_839 = s1_valid & T_833;
  assign T_840 = state == 2'h0;
  assign out_valid = T_839 & T_840;
  assign s1_idx = s1_vaddr[12:6];
  assign s1_hit = out_valid & s1_any_tag_hit;
  assign T_842 = s1_any_tag_hit == 1'h0;
  assign s1_miss = out_valid & T_842;
  assign T_845 = s1_miss == 1'h0;
  assign T_846 = T_840 & T_845;
  assign T_848 = s1_miss & T_840;
  assign GEN_1 = T_848 ? s1_paddr : refill_addr;
  assign refill_tag = refill_addr[31:13];
  assign FlowThroughSerializer_1_clk = clk;
  assign FlowThroughSerializer_1_reset = reset;
  assign FlowThroughSerializer_1_io_in_valid = io_mem_grant_valid;
  assign FlowThroughSerializer_1_io_in_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign FlowThroughSerializer_1_io_in_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign FlowThroughSerializer_1_io_in_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign FlowThroughSerializer_1_io_in_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign FlowThroughSerializer_1_io_in_bits_g_type = io_mem_grant_bits_g_type;
  assign FlowThroughSerializer_1_io_in_bits_data = io_mem_grant_bits_data;
  assign FlowThroughSerializer_1_io_out_ready = 1'h1;
  assign T_849 = FlowThroughSerializer_1_io_out_ready & FlowThroughSerializer_1_io_out_valid;
  assign T_852 = refill_cnt == 3'h7;
  assign T_854 = refill_cnt + 3'h1;
  assign T_855 = T_854[2:0];
  assign GEN_2 = T_849 ? T_855 : refill_cnt;
  assign refill_wrap = T_849 & T_852;
  assign T_856 = state == 2'h3;
  assign refill_done = T_856 & refill_wrap;
  assign tag_array_0_tag_rdata_addr = T_871;
  assign tag_array_0_tag_rdata_en = 1'h1;
  assign tag_array_0_tag_rdata_data = tag_array_0[GEN_11];
  assign tag_array_0_T_893_data = T_880_0;
  assign tag_array_0_T_893_addr = s1_idx;
  assign tag_array_0_T_893_mask = GEN_12;
  assign tag_array_0_T_893_en = refill_done;
  assign T_866 = s0_vaddr[12:6];
  assign T_871 = T_866;
  assign T_880_0 = refill_tag;
  assign T_889_0 = 1'h1;
  assign GEN_12 = refill_done ? T_889_0 : 1'h0;
  assign T_897 = invalidated == 1'h0;
  assign T_898 = refill_done & T_897;
  assign T_899 = {1'h0,s1_idx};
  assign T_902 = 256'h1 << T_899;
  assign GEN_36 = {{128'd0}, vb_array};
  assign T_903 = GEN_36 | T_902;
  assign T_904 = ~ vb_array;
  assign GEN_37 = {{128'd0}, T_904};
  assign T_905 = GEN_37 | T_902;
  assign T_906 = ~ T_905;
  assign GEN_13 = T_898 ? T_903 : {{128'd0}, vb_array};
  assign GEN_14 = io_invalidate ? 256'h0 : GEN_13;
  assign GEN_15 = io_invalidate ? 1'h1 : invalidated;
  assign s1_disparity_0 = 1'h0;
  assign T_917 = s1_valid & s1_disparity_0;
  assign GEN_16 = T_917 ? T_906 : GEN_14;
  assign s1_tag_match_0 = T_962;
  assign s1_tag_hit_0 = T_963;
  assign s1_dout_0 = T_974_T_987_data;
  assign T_950 = io_invalidate == 1'h0;
  assign T_954 = vb_array >> T_899;
  assign T_955 = T_954[0];
  assign T_957 = T_950 & T_955;
  assign T_961 = tag_array_0_tag_rdata_data;
  assign T_962 = T_961 == s1_tag;
  assign T_963 = T_957 & s1_tag_match_0;
  assign T_970 = s1_disparity_0 == 1'h0;
  assign T_971 = s1_tag_hit_0 & T_970;
  assign T_974_T_987_addr = T_986;
  assign T_974_T_987_en = 1'h1;
  assign T_974_T_987_data = T_974[GEN_38];
  assign T_974_T_980_data = GEN_20;
  assign T_974_T_980_addr = T_979;
  assign T_974_T_980_mask = T_977;
  assign T_974_T_980_en = T_977;
  assign T_977 = FlowThroughSerializer_1_io_out_valid;
  assign GEN_40 = {{3'd0}, s1_idx};
  assign T_978 = GEN_40 << 3;
  assign GEN_41 = {{7'd0}, refill_cnt};
  assign T_979 = T_978 | GEN_41;
  assign GEN_20 = FlowThroughSerializer_1_io_out_bits_data;
  assign T_981 = s0_vaddr[12:3];
  assign T_986 = T_981;
  assign T_989 = stall == 1'h0;
  assign GEN_23 = T_989 ? s1_hit : T_990;
  assign GEN_24 = T_989 ? s1_tag_hit_0 : T_995_0;
  assign GEN_25 = T_989 ? s1_dout_0 : T_1001_0;
  assign T_1003 = state == 2'h1;
  assign T_1005 = io_s2_kill == 1'h0;
  assign T_1006 = T_1003 & T_1005;
  assign T_1007 = refill_addr[31:6];
  assign T_1110_addr_block = T_1007;
  assign T_1110_client_xact_id = 1'h0;
  assign T_1110_addr_beat = 3'h0;
  assign T_1110_is_builtin_type = 1'h1;
  assign T_1110_a_type = 3'h1;
  assign T_1110_union = 12'h1c1;
  assign T_1110_data = 64'h0;
  assign T_1138 = 2'h0 == state;
  assign GEN_26 = s1_miss ? 2'h1 : state;
  assign GEN_27 = T_1138 ? GEN_26 : state;
  assign GEN_28 = T_1138 ? 1'h0 : GEN_15;
  assign T_1140 = 2'h1 == state;
  assign GEN_29 = io_mem_acquire_ready ? 2'h2 : GEN_27;
  assign GEN_30 = io_s2_kill ? 2'h0 : GEN_29;
  assign GEN_31 = T_1140 ? GEN_30 : GEN_27;
  assign T_1141 = 2'h2 == state;
  assign GEN_32 = io_mem_grant_valid ? 2'h3 : GEN_31;
  assign GEN_33 = T_1141 ? GEN_32 : GEN_31;
  assign T_1142 = 2'h3 == state;
  assign GEN_34 = refill_done ? 2'h0 : GEN_33;
  assign GEN_35 = T_1142 ? GEN_34 : GEN_33;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_4 = {1{$random}};
  state = GEN_4[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_5 = {1{$random}};
  invalidated = GEN_5[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_6 = {1{$random}};
  refill_addr = GEN_6[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_7 = {1{$random}};
  s1_valid = GEN_7[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_8 = {1{$random}};
  s1_vaddr = GEN_8[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_9 = {1{$random}};
  refill_cnt = GEN_9[2:0];
  `endif
  GEN_10 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tag_array_0[initvar] = GEN_10[18:0];
  `endif
  `ifdef RANDOMIZE
  GEN_17 = {1{$random}};
  GEN_11 = GEN_17[6:0];
  `endif
  `ifdef RANDOMIZE
  GEN_19 = {1{$random}};
  GEN_18 = GEN_19[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_21 = {4{$random}};
  vb_array = GEN_21[127:0];
  `endif
  GEN_22 = {2{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    T_974[initvar] = GEN_22[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_39 = {1{$random}};
  GEN_38 = GEN_39[9:0];
  `endif
  `ifdef RANDOMIZE
  GEN_43 = {1{$random}};
  GEN_42 = GEN_43[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_44 = {1{$random}};
  T_990 = GEN_44[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_45 = {1{$random}};
  T_995_0 = GEN_45[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_46 = {2{$random}};
  T_1001_0 = GEN_46[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_47 = {1{$random}};
  GEN_3 = GEN_47[31:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 2'h0;
    end else begin
      if(T_1142) begin
        if(refill_done) begin
          state <= 2'h0;
        end else begin
          if(T_1141) begin
            if(io_mem_grant_valid) begin
              state <= 2'h3;
            end else begin
              if(T_1140) begin
                if(io_s2_kill) begin
                  state <= 2'h0;
                end else begin
                  if(io_mem_acquire_ready) begin
                    state <= 2'h2;
                  end else begin
                    if(T_1138) begin
                      if(s1_miss) begin
                        state <= 2'h1;
                      end
                    end
                  end
                end
              end else begin
                if(T_1138) begin
                  if(s1_miss) begin
                    state <= 2'h1;
                  end
                end
              end
            end
          end else begin
            if(T_1140) begin
              if(io_s2_kill) begin
                state <= 2'h0;
              end else begin
                if(io_mem_acquire_ready) begin
                  state <= 2'h2;
                end else begin
                  if(T_1138) begin
                    if(s1_miss) begin
                      state <= 2'h1;
                    end
                  end
                end
              end
            end else begin
              if(T_1138) begin
                if(s1_miss) begin
                  state <= 2'h1;
                end
              end
            end
          end
        end
      end else begin
        if(T_1141) begin
          if(io_mem_grant_valid) begin
            state <= 2'h3;
          end else begin
            if(T_1140) begin
              if(io_s2_kill) begin
                state <= 2'h0;
              end else begin
                if(io_mem_acquire_ready) begin
                  state <= 2'h2;
                end else begin
                  state <= GEN_27;
                end
              end
            end else begin
              state <= GEN_27;
            end
          end
        end else begin
          if(T_1140) begin
            if(io_s2_kill) begin
              state <= 2'h0;
            end else begin
              if(io_mem_acquire_ready) begin
                state <= 2'h2;
              end else begin
                state <= GEN_27;
              end
            end
          end else begin
            state <= GEN_27;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1138) begin
        invalidated <= 1'h0;
      end else begin
        if(io_invalidate) begin
          invalidated <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_848) begin
        refill_addr <= s1_paddr;
      end
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T_835;
    end
    if(1'h0) begin
    end else begin
      if(T_830) begin
        s1_vaddr <= io_req_bits_addr;
      end
    end
    if(reset) begin
      refill_cnt <= 3'h0;
    end else begin
      if(T_849) begin
        refill_cnt <= T_855;
      end
    end
    GEN_11 <= tag_array_0_tag_rdata_addr;
    GEN_18 <= tag_array_0_tag_rdata_en;
    if(tag_array_0_T_893_en & tag_array_0_T_893_mask) begin
      tag_array_0[tag_array_0_T_893_addr] <= tag_array_0_T_893_data;
    end
    if(reset) begin
      vb_array <= 128'h0;
    end else begin
      vb_array <= GEN_16[127:0];
    end
    GEN_38 <= T_974_T_987_addr;
    GEN_42 <= T_974_T_987_en;
    if(T_974_T_980_en & T_974_T_980_mask) begin
      T_974[T_974_T_980_addr] <= T_974_T_980_data;
    end
    if(1'h0) begin
    end else begin
      if(T_989) begin
        T_990 <= s1_hit;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_989) begin
        T_995_0 <= s1_tag_hit_0;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_989) begin
        T_1001_0 <= s1_dout_0;
      end
    end
  end
endmodule
module TLB(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [19:0] io_req_bits_vpn,
  input   io_req_bits_passthrough,
  input   io_req_bits_instruction,
  input   io_req_bits_store,
  output  io_resp_miss,
  output [19:0] io_resp_ppn,
  output  io_resp_xcpt_ld,
  output  io_resp_xcpt_st,
  output  io_resp_xcpt_if,
  output  io_resp_cacheable,
  input   io_ptw_req_ready,
  output  io_ptw_req_valid,
  output [1:0] io_ptw_req_bits_prv,
  output  io_ptw_req_bits_pum,
  output  io_ptw_req_bits_mxr,
  output [19:0] io_ptw_req_bits_addr,
  output  io_ptw_req_bits_store,
  output  io_ptw_req_bits_fetch,
  input   io_ptw_resp_valid,
  input  [15:0] io_ptw_resp_bits_pte_reserved_for_hardware,
  input  [37:0] io_ptw_resp_bits_pte_ppn,
  input  [1:0] io_ptw_resp_bits_pte_reserved_for_software,
  input   io_ptw_resp_bits_pte_d,
  input   io_ptw_resp_bits_pte_a,
  input   io_ptw_resp_bits_pte_g,
  input   io_ptw_resp_bits_pte_u,
  input   io_ptw_resp_bits_pte_x,
  input   io_ptw_resp_bits_pte_w,
  input   io_ptw_resp_bits_pte_r,
  input   io_ptw_resp_bits_pte_v,
  input  [6:0] io_ptw_ptbr_asid,
  input  [21:0] io_ptw_ptbr_ppn,
  input   io_ptw_invalidate,
  input   io_ptw_status_debug,
  input  [1:0] io_ptw_status_prv,
  input   io_ptw_status_sd,
  input  [30:0] io_ptw_status_zero3,
  input   io_ptw_status_sd_rv32,
  input  [1:0] io_ptw_status_zero2,
  input  [4:0] io_ptw_status_vm,
  input  [3:0] io_ptw_status_zero1,
  input   io_ptw_status_mxr,
  input   io_ptw_status_pum,
  input   io_ptw_status_mprv,
  input  [1:0] io_ptw_status_xs,
  input  [1:0] io_ptw_status_fs,
  input  [1:0] io_ptw_status_mpp,
  input  [1:0] io_ptw_status_hpp,
  input   io_ptw_status_spp,
  input   io_ptw_status_mpie,
  input   io_ptw_status_hpie,
  input   io_ptw_status_spie,
  input   io_ptw_status_upie,
  input   io_ptw_status_mie,
  input   io_ptw_status_hie,
  input   io_ptw_status_sie,
  input   io_ptw_status_uie
);
  reg [3:0] valid;
  reg [31:0] GEN_10;
  reg [37:0] ppns_0;
  reg [63:0] GEN_15;
  reg [37:0] ppns_1;
  reg [63:0] GEN_26;
  reg [37:0] ppns_2;
  reg [63:0] GEN_27;
  reg [37:0] ppns_3;
  reg [63:0] GEN_28;
  reg [26:0] tags_0;
  reg [31:0] GEN_29;
  reg [26:0] tags_1;
  reg [31:0] GEN_30;
  reg [26:0] tags_2;
  reg [31:0] GEN_31;
  reg [26:0] tags_3;
  reg [31:0] GEN_32;
  reg [1:0] state;
  reg [31:0] GEN_33;
  reg [26:0] r_refill_tag;
  reg [31:0] GEN_34;
  reg [1:0] r_refill_waddr;
  reg [31:0] GEN_35;
  reg [19:0] r_req_vpn;
  reg [31:0] GEN_36;
  reg  r_req_passthrough;
  reg [31:0] GEN_37;
  reg  r_req_instruction;
  reg [31:0] GEN_38;
  reg  r_req_store;
  reg [31:0] GEN_39;
  wire [26:0] lookup_tag;
  wire  T_216;
  wire  T_217;
  wire  T_218;
  wire  T_219;
  wire  T_220;
  wire  T_221;
  wire  T_222;
  wire  T_223;
  wire  T_224;
  wire  T_225;
  wire  T_226;
  wire  T_227;
  reg [15:0] pte_array_reserved_for_hardware;
  reg [31:0] GEN_40;
  reg [37:0] pte_array_ppn;
  reg [63:0] GEN_41;
  reg [1:0] pte_array_reserved_for_software;
  reg [31:0] GEN_42;
  reg  pte_array_d;
  reg [31:0] GEN_43;
  reg  pte_array_a;
  reg [31:0] GEN_44;
  reg  pte_array_g;
  reg [31:0] GEN_45;
  reg  pte_array_u;
  reg [31:0] GEN_46;
  reg  pte_array_x;
  reg [31:0] GEN_47;
  reg  pte_array_w;
  reg [31:0] GEN_48;
  reg  pte_array_r;
  reg [31:0] GEN_49;
  reg  pte_array_v;
  reg [31:0] GEN_50;
  reg [3:0] u_array;
  reg [31:0] GEN_51;
  reg [3:0] sw_array;
  reg [31:0] GEN_52;
  reg [3:0] sx_array;
  reg [31:0] GEN_53;
  reg [3:0] sr_array;
  reg [31:0] GEN_54;
  reg [3:0] dirty_array;
  reg [31:0] GEN_55;
  wire [37:0] GEN_0;
  wire [37:0] GEN_2;
  wire [37:0] GEN_3;
  wire [37:0] GEN_4;
  wire [37:0] GEN_5;
  wire [26:0] GEN_1;
  wire [26:0] GEN_6;
  wire [26:0] GEN_7;
  wire [26:0] GEN_8;
  wire [26:0] GEN_9;
  wire [3:0] T_259;
  wire [3:0] T_260;
  wire [3:0] T_261;
  wire [3:0] T_262;
  wire [3:0] T_263;
  wire [3:0] T_264;
  wire  T_266;
  wire  T_267;
  wire  T_268;
  wire  T_269;
  wire  T_270;
  wire [3:0] T_271;
  wire [3:0] T_273;
  wire [3:0] T_274;
  wire  T_280;
  wire [3:0] T_281;
  wire [3:0] T_283;
  wire [3:0] T_284;
  wire  T_290;
  wire [3:0] T_291;
  wire [3:0] T_293;
  wire [3:0] T_294;
  wire [3:0] T_295;
  wire [3:0] T_297;
  wire [3:0] T_298;
  wire [37:0] GEN_11;
  wire [37:0] GEN_12;
  wire [37:0] GEN_13;
  wire [37:0] GEN_14;
  wire [26:0] GEN_16;
  wire [26:0] GEN_17;
  wire [26:0] GEN_18;
  wire [26:0] GEN_19;
  wire [3:0] GEN_20;
  wire [3:0] GEN_21;
  wire [3:0] GEN_22;
  wire [3:0] GEN_23;
  wire [3:0] GEN_24;
  wire [3:0] GEN_25;
  reg [3:0] T_300;
  reg [31:0] GEN_56;
  wire [31:0] paddr;
  wire  T_390;
  wire [2:0] T_394;
  wire  T_396;
  wire  T_398;
  wire  T_399;
  wire [2:0] T_402;
  wire  T_404;
  wire  T_406;
  wire  T_407;
  wire [2:0] T_410;
  wire  T_412;
  wire  T_414;
  wire  T_415;
  wire [2:0] T_418;
  wire  T_420;
  wire  T_422;
  wire  T_423;
  wire [2:0] T_426;
  wire  T_428;
  wire  T_430;
  wire  T_431;
  wire [2:0] T_434;
  wire [2:0] T_439;
  wire [2:0] T_440;
  wire [2:0] T_441;
  wire [2:0] T_442;
  wire [2:0] T_443;
  wire  addr_prot_x;
  wire  addr_prot_w;
  wire  addr_prot_r;
  wire  T_451;
  wire  T_452;
  wire  T_453;
  wire  T_454;
  wire  T_458;
  wire  T_471;
  wire  T_484;
  wire [37:0] T_502;
  wire [37:0] T_504;
  wire [37:0] T_506;
  wire [37:0] T_508;
  wire [37:0] T_510;
  wire [37:0] T_511;
  wire [37:0] T_512;
  wire [37:0] T_513;
  wire [37:0] T_515;
  wire  T_516;
  assign io_req_ready = T_454;
  assign io_resp_miss = 1'h0;
  assign io_resp_ppn = T_515[19:0];
  assign io_resp_xcpt_ld = T_458;
  assign io_resp_xcpt_st = T_471;
  assign io_resp_xcpt_if = T_484;
  assign io_resp_cacheable = T_431;
  assign io_ptw_req_valid = T_516;
  assign io_ptw_req_bits_prv = io_ptw_status_prv;
  assign io_ptw_req_bits_pum = io_ptw_status_pum;
  assign io_ptw_req_bits_mxr = io_ptw_status_mxr;
  assign io_ptw_req_bits_addr = r_refill_tag[19:0];
  assign io_ptw_req_bits_store = r_req_store;
  assign io_ptw_req_bits_fetch = r_req_instruction;
  assign lookup_tag = {io_ptw_ptbr_asid,io_req_bits_vpn};
  assign T_216 = valid[0];
  assign T_217 = tags_0 == lookup_tag;
  assign T_218 = T_216 & T_217;
  assign T_219 = valid[1];
  assign T_220 = tags_1 == lookup_tag;
  assign T_221 = T_219 & T_220;
  assign T_222 = valid[2];
  assign T_223 = tags_2 == lookup_tag;
  assign T_224 = T_222 & T_223;
  assign T_225 = valid[3];
  assign T_226 = tags_3 == lookup_tag;
  assign T_227 = T_225 & T_226;
  assign GEN_0 = io_ptw_resp_bits_pte_ppn;
  assign GEN_2 = 2'h0 == r_refill_waddr ? GEN_0 : ppns_0;
  assign GEN_3 = 2'h1 == r_refill_waddr ? GEN_0 : ppns_1;
  assign GEN_4 = 2'h2 == r_refill_waddr ? GEN_0 : ppns_2;
  assign GEN_5 = 2'h3 == r_refill_waddr ? GEN_0 : ppns_3;
  assign GEN_1 = r_refill_tag;
  assign GEN_6 = 2'h0 == r_refill_waddr ? GEN_1 : tags_0;
  assign GEN_7 = 2'h1 == r_refill_waddr ? GEN_1 : tags_1;
  assign GEN_8 = 2'h2 == r_refill_waddr ? GEN_1 : tags_2;
  assign GEN_9 = 2'h3 == r_refill_waddr ? GEN_1 : tags_3;
  assign T_259 = 4'h1 << r_refill_waddr;
  assign T_260 = valid | T_259;
  assign T_261 = u_array | T_259;
  assign T_262 = ~ T_259;
  assign T_263 = u_array & T_262;
  assign T_264 = io_ptw_resp_bits_pte_u ? T_261 : T_263;
  assign T_266 = io_ptw_resp_bits_pte_w == 1'h0;
  assign T_267 = io_ptw_resp_bits_pte_x & T_266;
  assign T_268 = io_ptw_resp_bits_pte_r | T_267;
  assign T_269 = io_ptw_resp_bits_pte_v & T_268;
  assign T_270 = T_269 & io_ptw_resp_bits_pte_r;
  assign T_271 = sr_array | T_259;
  assign T_273 = sr_array & T_262;
  assign T_274 = T_270 ? T_271 : T_273;
  assign T_280 = T_269 & io_ptw_resp_bits_pte_w;
  assign T_281 = sw_array | T_259;
  assign T_283 = sw_array & T_262;
  assign T_284 = T_280 ? T_281 : T_283;
  assign T_290 = T_269 & io_ptw_resp_bits_pte_x;
  assign T_291 = sx_array | T_259;
  assign T_293 = sx_array & T_262;
  assign T_294 = T_290 ? T_291 : T_293;
  assign T_295 = dirty_array | T_259;
  assign T_297 = dirty_array & T_262;
  assign T_298 = io_ptw_resp_bits_pte_d ? T_295 : T_297;
  assign GEN_11 = io_ptw_resp_valid ? GEN_2 : ppns_0;
  assign GEN_12 = io_ptw_resp_valid ? GEN_3 : ppns_1;
  assign GEN_13 = io_ptw_resp_valid ? GEN_4 : ppns_2;
  assign GEN_14 = io_ptw_resp_valid ? GEN_5 : ppns_3;
  assign GEN_16 = io_ptw_resp_valid ? GEN_6 : tags_0;
  assign GEN_17 = io_ptw_resp_valid ? GEN_7 : tags_1;
  assign GEN_18 = io_ptw_resp_valid ? GEN_8 : tags_2;
  assign GEN_19 = io_ptw_resp_valid ? GEN_9 : tags_3;
  assign GEN_20 = io_ptw_resp_valid ? T_260 : valid;
  assign GEN_21 = io_ptw_resp_valid ? T_264 : u_array;
  assign GEN_22 = io_ptw_resp_valid ? T_274 : sr_array;
  assign GEN_23 = io_ptw_resp_valid ? T_284 : sw_array;
  assign GEN_24 = io_ptw_resp_valid ? T_294 : sx_array;
  assign GEN_25 = io_ptw_resp_valid ? T_298 : dirty_array;
  assign paddr = {io_resp_ppn,12'h0};
  assign T_390 = paddr < 32'h1000;
  assign T_394 = T_390 ? 3'h7 : 3'h0;
  assign T_396 = 32'h1000 <= paddr;
  assign T_398 = paddr < 32'h2000;
  assign T_399 = T_396 & T_398;
  assign T_402 = T_399 ? 3'h5 : 3'h0;
  assign T_404 = 32'h40000000 <= paddr;
  assign T_406 = paddr < 32'h44000000;
  assign T_407 = T_404 & T_406;
  assign T_410 = T_407 ? 3'h3 : 3'h0;
  assign T_412 = 32'h44000000 <= paddr;
  assign T_414 = paddr < 32'h48000000;
  assign T_415 = T_412 & T_414;
  assign T_418 = T_415 ? 3'h3 : 3'h0;
  assign T_420 = 32'h60000000 <= paddr;
  assign T_422 = paddr < 32'h80000000;
  assign T_423 = T_420 & T_422;
  assign T_426 = T_423 ? 3'h7 : 3'h0;
  assign T_428 = 32'h80000000 <= paddr;
  assign T_430 = paddr < 32'h90000000;
  assign T_431 = T_428 & T_430;
  assign T_434 = T_431 ? 3'h7 : 3'h0;
  assign T_439 = T_394 | T_402;
  assign T_440 = T_439 | T_410;
  assign T_441 = T_440 | T_418;
  assign T_442 = T_441 | T_426;
  assign T_443 = T_442 | T_434;
  assign addr_prot_x = T_453;
  assign addr_prot_w = T_452;
  assign addr_prot_r = T_451;
  assign T_451 = T_443[0];
  assign T_452 = T_443[1];
  assign T_453 = T_443[2];
  assign T_454 = state == 2'h0;
  assign T_458 = addr_prot_r == 1'h0;
  assign T_471 = addr_prot_w == 1'h0;
  assign T_484 = addr_prot_x == 1'h0;
  assign T_502 = T_218 ? ppns_0 : 38'h0;
  assign T_504 = T_221 ? ppns_1 : 38'h0;
  assign T_506 = T_224 ? ppns_2 : 38'h0;
  assign T_508 = T_227 ? ppns_3 : 38'h0;
  assign T_510 = T_502 | T_504;
  assign T_511 = T_510 | T_506;
  assign T_512 = T_511 | T_508;
  assign T_513 = T_512;
  assign T_515 = {{18'd0}, io_req_bits_vpn};
  assign T_516 = state == 2'h1;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_10 = {1{$random}};
  valid = GEN_10[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_15 = {2{$random}};
  ppns_0 = GEN_15[37:0];
  `endif
  `ifdef RANDOMIZE
  GEN_26 = {2{$random}};
  ppns_1 = GEN_26[37:0];
  `endif
  `ifdef RANDOMIZE
  GEN_27 = {2{$random}};
  ppns_2 = GEN_27[37:0];
  `endif
  `ifdef RANDOMIZE
  GEN_28 = {2{$random}};
  ppns_3 = GEN_28[37:0];
  `endif
  `ifdef RANDOMIZE
  GEN_29 = {1{$random}};
  tags_0 = GEN_29[26:0];
  `endif
  `ifdef RANDOMIZE
  GEN_30 = {1{$random}};
  tags_1 = GEN_30[26:0];
  `endif
  `ifdef RANDOMIZE
  GEN_31 = {1{$random}};
  tags_2 = GEN_31[26:0];
  `endif
  `ifdef RANDOMIZE
  GEN_32 = {1{$random}};
  tags_3 = GEN_32[26:0];
  `endif
  `ifdef RANDOMIZE
  GEN_33 = {1{$random}};
  state = GEN_33[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_34 = {1{$random}};
  r_refill_tag = GEN_34[26:0];
  `endif
  `ifdef RANDOMIZE
  GEN_35 = {1{$random}};
  r_refill_waddr = GEN_35[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_36 = {1{$random}};
  r_req_vpn = GEN_36[19:0];
  `endif
  `ifdef RANDOMIZE
  GEN_37 = {1{$random}};
  r_req_passthrough = GEN_37[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_38 = {1{$random}};
  r_req_instruction = GEN_38[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_39 = {1{$random}};
  r_req_store = GEN_39[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_40 = {1{$random}};
  pte_array_reserved_for_hardware = GEN_40[15:0];
  `endif
  `ifdef RANDOMIZE
  GEN_41 = {2{$random}};
  pte_array_ppn = GEN_41[37:0];
  `endif
  `ifdef RANDOMIZE
  GEN_42 = {1{$random}};
  pte_array_reserved_for_software = GEN_42[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_43 = {1{$random}};
  pte_array_d = GEN_43[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_44 = {1{$random}};
  pte_array_a = GEN_44[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_45 = {1{$random}};
  pte_array_g = GEN_45[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_46 = {1{$random}};
  pte_array_u = GEN_46[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_47 = {1{$random}};
  pte_array_x = GEN_47[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_48 = {1{$random}};
  pte_array_w = GEN_48[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_49 = {1{$random}};
  pte_array_r = GEN_49[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_50 = {1{$random}};
  pte_array_v = GEN_50[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_51 = {1{$random}};
  u_array = GEN_51[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_52 = {1{$random}};
  sw_array = GEN_52[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_53 = {1{$random}};
  sx_array = GEN_53[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_54 = {1{$random}};
  sr_array = GEN_54[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_55 = {1{$random}};
  dirty_array = GEN_55[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_56 = {1{$random}};
  T_300 = GEN_56[3:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      valid <= 4'h0;
    end else begin
      if(io_ptw_resp_valid) begin
        valid <= T_260;
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(2'h0 == r_refill_waddr) begin
          ppns_0 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(2'h1 == r_refill_waddr) begin
          ppns_1 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(2'h2 == r_refill_waddr) begin
          ppns_2 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(2'h3 == r_refill_waddr) begin
          ppns_3 <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(2'h0 == r_refill_waddr) begin
          tags_0 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(2'h1 == r_refill_waddr) begin
          tags_1 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(2'h2 == r_refill_waddr) begin
          tags_2 <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(2'h3 == r_refill_waddr) begin
          tags_3 <= GEN_1;
        end
      end
    end
    if(reset) begin
      state <= 2'h0;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(io_ptw_resp_bits_pte_u) begin
          u_array <= T_261;
        end else begin
          u_array <= T_263;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(T_280) begin
          sw_array <= T_281;
        end else begin
          sw_array <= T_283;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(T_290) begin
          sx_array <= T_291;
        end else begin
          sx_array <= T_293;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(T_270) begin
          sr_array <= T_271;
        end else begin
          sr_array <= T_273;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_ptw_resp_valid) begin
        if(io_ptw_resp_bits_pte_d) begin
          dirty_array <= T_295;
        end else begin
          dirty_array <= T_297;
        end
      end
    end
    if(1'h0) begin
    end
  end
endmodule
module Frontend(
  input   clk,
  input   reset,
  input   io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_pc,
  input   io_cpu_req_bits_speculative,
  input   io_cpu_resp_ready,
  output  io_cpu_resp_valid,
  output [31:0] io_cpu_resp_bits_pc,
  output [31:0] io_cpu_resp_bits_data_0,
  output  io_cpu_resp_bits_mask,
  output  io_cpu_resp_bits_xcpt_if,
  output  io_cpu_resp_bits_replay,
  output  io_cpu_btb_resp_valid,
  output  io_cpu_btb_resp_bits_taken,
  output  io_cpu_btb_resp_bits_mask,
  output  io_cpu_btb_resp_bits_bridx,
  output [31:0] io_cpu_btb_resp_bits_target,
  output  io_cpu_btb_resp_bits_entry,
  output  io_cpu_btb_resp_bits_bht_history,
  output [1:0] io_cpu_btb_resp_bits_bht_value,
  input   io_cpu_btb_update_valid,
  input   io_cpu_btb_update_bits_prediction_valid,
  input   io_cpu_btb_update_bits_prediction_bits_taken,
  input   io_cpu_btb_update_bits_prediction_bits_mask,
  input   io_cpu_btb_update_bits_prediction_bits_bridx,
  input  [31:0] io_cpu_btb_update_bits_prediction_bits_target,
  input   io_cpu_btb_update_bits_prediction_bits_entry,
  input   io_cpu_btb_update_bits_prediction_bits_bht_history,
  input  [1:0] io_cpu_btb_update_bits_prediction_bits_bht_value,
  input  [31:0] io_cpu_btb_update_bits_pc,
  input  [31:0] io_cpu_btb_update_bits_target,
  input   io_cpu_btb_update_bits_taken,
  input   io_cpu_btb_update_bits_isJump,
  input   io_cpu_btb_update_bits_isReturn,
  input  [31:0] io_cpu_btb_update_bits_br_pc,
  input   io_cpu_bht_update_valid,
  input   io_cpu_bht_update_bits_prediction_valid,
  input   io_cpu_bht_update_bits_prediction_bits_taken,
  input   io_cpu_bht_update_bits_prediction_bits_mask,
  input   io_cpu_bht_update_bits_prediction_bits_bridx,
  input  [31:0] io_cpu_bht_update_bits_prediction_bits_target,
  input   io_cpu_bht_update_bits_prediction_bits_entry,
  input   io_cpu_bht_update_bits_prediction_bits_bht_history,
  input  [1:0] io_cpu_bht_update_bits_prediction_bits_bht_value,
  input  [31:0] io_cpu_bht_update_bits_pc,
  input   io_cpu_bht_update_bits_taken,
  input   io_cpu_bht_update_bits_mispredict,
  input   io_cpu_ras_update_valid,
  input   io_cpu_ras_update_bits_isCall,
  input   io_cpu_ras_update_bits_isReturn,
  input  [31:0] io_cpu_ras_update_bits_returnAddr,
  input   io_cpu_ras_update_bits_prediction_valid,
  input   io_cpu_ras_update_bits_prediction_bits_taken,
  input   io_cpu_ras_update_bits_prediction_bits_mask,
  input   io_cpu_ras_update_bits_prediction_bits_bridx,
  input  [31:0] io_cpu_ras_update_bits_prediction_bits_target,
  input   io_cpu_ras_update_bits_prediction_bits_entry,
  input   io_cpu_ras_update_bits_prediction_bits_bht_history,
  input  [1:0] io_cpu_ras_update_bits_prediction_bits_bht_value,
  input   io_cpu_flush_icache,
  input   io_cpu_flush_tlb,
  output [31:0] io_cpu_npc,
  input   io_ptw_req_ready,
  output  io_ptw_req_valid,
  output [1:0] io_ptw_req_bits_prv,
  output  io_ptw_req_bits_pum,
  output  io_ptw_req_bits_mxr,
  output [19:0] io_ptw_req_bits_addr,
  output  io_ptw_req_bits_store,
  output  io_ptw_req_bits_fetch,
  input   io_ptw_resp_valid,
  input  [15:0] io_ptw_resp_bits_pte_reserved_for_hardware,
  input  [37:0] io_ptw_resp_bits_pte_ppn,
  input  [1:0] io_ptw_resp_bits_pte_reserved_for_software,
  input   io_ptw_resp_bits_pte_d,
  input   io_ptw_resp_bits_pte_a,
  input   io_ptw_resp_bits_pte_g,
  input   io_ptw_resp_bits_pte_u,
  input   io_ptw_resp_bits_pte_x,
  input   io_ptw_resp_bits_pte_w,
  input   io_ptw_resp_bits_pte_r,
  input   io_ptw_resp_bits_pte_v,
  input  [6:0] io_ptw_ptbr_asid,
  input  [21:0] io_ptw_ptbr_ppn,
  input   io_ptw_invalidate,
  input   io_ptw_status_debug,
  input  [1:0] io_ptw_status_prv,
  input   io_ptw_status_sd,
  input  [30:0] io_ptw_status_zero3,
  input   io_ptw_status_sd_rv32,
  input  [1:0] io_ptw_status_zero2,
  input  [4:0] io_ptw_status_vm,
  input  [3:0] io_ptw_status_zero1,
  input   io_ptw_status_mxr,
  input   io_ptw_status_pum,
  input   io_ptw_status_mprv,
  input  [1:0] io_ptw_status_xs,
  input  [1:0] io_ptw_status_fs,
  input  [1:0] io_ptw_status_mpp,
  input  [1:0] io_ptw_status_hpp,
  input   io_ptw_status_spp,
  input   io_ptw_status_mpie,
  input   io_ptw_status_hpie,
  input   io_ptw_status_spie,
  input   io_ptw_status_upie,
  input   io_ptw_status_mie,
  input   io_ptw_status_hie,
  input   io_ptw_status_sie,
  input   io_ptw_status_uie,
  input   io_mem_acquire_ready,
  output  io_mem_acquire_valid,
  output [25:0] io_mem_acquire_bits_addr_block,
  output  io_mem_acquire_bits_client_xact_id,
  output [2:0] io_mem_acquire_bits_addr_beat,
  output  io_mem_acquire_bits_is_builtin_type,
  output [2:0] io_mem_acquire_bits_a_type,
  output [11:0] io_mem_acquire_bits_union,
  output [63:0] io_mem_acquire_bits_data,
  output  io_mem_grant_ready,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input   io_mem_grant_bits_client_xact_id,
  input  [1:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data
);
//<CJ> RESET_VECTOR_ADDR
  parameter RESET_VECTOR_ADDR = 60000000;

  wire  icache_clk;
  wire  icache_reset;
  wire  icache_io_req_valid;
  wire [31:0] icache_io_req_bits_addr;
  wire [19:0] icache_io_s1_ppn;
  wire  icache_io_s1_kill;
  wire  icache_io_s2_kill;
  wire  icache_io_resp_ready;
  wire  icache_io_resp_valid;
  wire [31:0] icache_io_resp_bits_data;
  wire [63:0] icache_io_resp_bits_datablock;
  wire  icache_io_invalidate;
  wire  icache_io_mem_acquire_ready;
  wire  icache_io_mem_acquire_valid;
  wire [25:0] icache_io_mem_acquire_bits_addr_block;
  wire  icache_io_mem_acquire_bits_client_xact_id;
  wire [2:0] icache_io_mem_acquire_bits_addr_beat;
  wire  icache_io_mem_acquire_bits_is_builtin_type;
  wire [2:0] icache_io_mem_acquire_bits_a_type;
  wire [11:0] icache_io_mem_acquire_bits_union;
  wire [63:0] icache_io_mem_acquire_bits_data;
  wire  icache_io_mem_grant_ready;
  wire  icache_io_mem_grant_valid;
  wire [2:0] icache_io_mem_grant_bits_addr_beat;
  wire  icache_io_mem_grant_bits_client_xact_id;
  wire [1:0] icache_io_mem_grant_bits_manager_xact_id;
  wire  icache_io_mem_grant_bits_is_builtin_type;
  wire [3:0] icache_io_mem_grant_bits_g_type;
  wire [63:0] icache_io_mem_grant_bits_data;
  wire  tlb_clk;
  wire  tlb_reset;
  wire  tlb_io_req_ready;
  wire  tlb_io_req_valid;
  wire [19:0] tlb_io_req_bits_vpn;
  wire  tlb_io_req_bits_passthrough;
  wire  tlb_io_req_bits_instruction;
  wire  tlb_io_req_bits_store;
  wire  tlb_io_resp_miss;
  wire [19:0] tlb_io_resp_ppn;
  wire  tlb_io_resp_xcpt_ld;
  wire  tlb_io_resp_xcpt_st;
  wire  tlb_io_resp_xcpt_if;
  wire  tlb_io_resp_cacheable;
  wire  tlb_io_ptw_req_ready;
  wire  tlb_io_ptw_req_valid;
  wire [1:0] tlb_io_ptw_req_bits_prv;
  wire  tlb_io_ptw_req_bits_pum;
  wire  tlb_io_ptw_req_bits_mxr;
  wire [19:0] tlb_io_ptw_req_bits_addr;
  wire  tlb_io_ptw_req_bits_store;
  wire  tlb_io_ptw_req_bits_fetch;
  wire  tlb_io_ptw_resp_valid;
  wire [15:0] tlb_io_ptw_resp_bits_pte_reserved_for_hardware;
  wire [37:0] tlb_io_ptw_resp_bits_pte_ppn;
  wire [1:0] tlb_io_ptw_resp_bits_pte_reserved_for_software;
  wire  tlb_io_ptw_resp_bits_pte_d;
  wire  tlb_io_ptw_resp_bits_pte_a;
  wire  tlb_io_ptw_resp_bits_pte_g;
  wire  tlb_io_ptw_resp_bits_pte_u;
  wire  tlb_io_ptw_resp_bits_pte_x;
  wire  tlb_io_ptw_resp_bits_pte_w;
  wire  tlb_io_ptw_resp_bits_pte_r;
  wire  tlb_io_ptw_resp_bits_pte_v;
  wire [6:0] tlb_io_ptw_ptbr_asid;
  wire [21:0] tlb_io_ptw_ptbr_ppn;
  wire  tlb_io_ptw_invalidate;
  wire  tlb_io_ptw_status_debug;
  wire [1:0] tlb_io_ptw_status_prv;
  wire  tlb_io_ptw_status_sd;
  wire [30:0] tlb_io_ptw_status_zero3;
  wire  tlb_io_ptw_status_sd_rv32;
  wire [1:0] tlb_io_ptw_status_zero2;
  wire [4:0] tlb_io_ptw_status_vm;
  wire [3:0] tlb_io_ptw_status_zero1;
  wire  tlb_io_ptw_status_mxr;
  wire  tlb_io_ptw_status_pum;
  wire  tlb_io_ptw_status_mprv;
  wire [1:0] tlb_io_ptw_status_xs;
  wire [1:0] tlb_io_ptw_status_fs;
  wire [1:0] tlb_io_ptw_status_mpp;
  wire [1:0] tlb_io_ptw_status_hpp;
  wire  tlb_io_ptw_status_spp;
  wire  tlb_io_ptw_status_mpie;
  wire  tlb_io_ptw_status_hpie;
  wire  tlb_io_ptw_status_spie;
  wire  tlb_io_ptw_status_upie;
  wire  tlb_io_ptw_status_mie;
  wire  tlb_io_ptw_status_hie;
  wire  tlb_io_ptw_status_sie;
  wire  tlb_io_ptw_status_uie;
  reg [31:0] s1_pc_;
  reg [31:0] GEN_15;
  wire [31:0] T_1315;
  wire [31:0] T_1317;
  wire [31:0] s1_pc;
  reg  s1_speculative;
  reg [31:0] GEN_16;
  reg  s1_same_block;
  reg [31:0] GEN_17;
  reg  s2_valid;
  reg [31:0] GEN_18;
  reg [31:0] s2_pc;
  reg [31:0] GEN_19;
  reg  s2_btb_resp_valid;
  reg [31:0] GEN_20;
  reg  s2_btb_resp_bits_taken;
  reg [31:0] GEN_21;
  reg  s2_btb_resp_bits_mask;
  reg [31:0] GEN_22;
  reg  s2_btb_resp_bits_bridx;
  reg [31:0] GEN_23;
  reg [31:0] s2_btb_resp_bits_target;
  reg [31:0] GEN_24;
  reg  s2_btb_resp_bits_entry;
  reg [31:0] GEN_25;
  reg  s2_btb_resp_bits_bht_history;
  reg [31:0] GEN_26;
  reg [1:0] s2_btb_resp_bits_bht_value;
  reg [31:0] GEN_27;
  reg  s2_xcpt_if;
  reg [31:0] GEN_28;
  reg  s2_speculative;
  reg [31:0] GEN_29;
  wire [31:0] T_1342;
  wire [31:0] T_1344;
  wire [31:0] T_1345;
  wire [32:0] T_1347;
  wire [31:0] ntpc;
  wire [31:0] predicted_npc;
  wire  T_1349;
  wire  icmiss;
  wire [31:0] npc;
  wire  T_1351;
  wire  T_1353;
  wire  T_1354;
  wire [31:0] T_1356;
  wire [31:0] T_1358;
  wire  T_1359;
  wire  T_1360;
  wire  s0_same_block;
  wire  T_1362;
  wire  stall;
  wire  T_1364;
  wire  T_1366;
  wire  T_1367;
  wire  T_1369;
  wire  T_1375;
  wire  T_1376;
  wire [31:0] GEN_0;
  wire  GEN_1;
  wire  GEN_2;
  wire  GEN_3;
  wire [31:0] GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire [31:0] GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire [31:0] GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  T_1383;
  wire [19:0] T_1384;
  wire  T_1391;
  wire  T_1392;
  wire  T_1393;
  wire  T_1394;
  wire  T_1395;
  wire  T_1396;
  wire  T_1400;
  wire  T_1401;
  wire  T_1402;
  wire  T_1403;
  wire  T_1404;
  wire [31:0] T_1405;
  wire  T_1406;
  wire [5:0] GEN_14;
  wire [5:0] T_1407;
  wire [63:0] fetch_data;
  wire [31:0] T_1408;
  wire [1:0] T_1411;
  wire  T_1414;
  wire  T_1416;
  wire  T_1417;
  ICache icache (
    .clk(icache_clk),
    .reset(icache_reset),
    .io_req_valid(icache_io_req_valid),
    .io_req_bits_addr(icache_io_req_bits_addr),
    .io_s1_ppn(icache_io_s1_ppn),
    .io_s1_kill(icache_io_s1_kill),
    .io_s2_kill(icache_io_s2_kill),
    .io_resp_ready(icache_io_resp_ready),
    .io_resp_valid(icache_io_resp_valid),
    .io_resp_bits_data(icache_io_resp_bits_data),
    .io_resp_bits_datablock(icache_io_resp_bits_datablock),
    .io_invalidate(icache_io_invalidate),
    .io_mem_acquire_ready(icache_io_mem_acquire_ready),
    .io_mem_acquire_valid(icache_io_mem_acquire_valid),
    .io_mem_acquire_bits_addr_block(icache_io_mem_acquire_bits_addr_block),
    .io_mem_acquire_bits_client_xact_id(icache_io_mem_acquire_bits_client_xact_id),
    .io_mem_acquire_bits_addr_beat(icache_io_mem_acquire_bits_addr_beat),
    .io_mem_acquire_bits_is_builtin_type(icache_io_mem_acquire_bits_is_builtin_type),
    .io_mem_acquire_bits_a_type(icache_io_mem_acquire_bits_a_type),
    .io_mem_acquire_bits_union(icache_io_mem_acquire_bits_union),
    .io_mem_acquire_bits_data(icache_io_mem_acquire_bits_data),
    .io_mem_grant_ready(icache_io_mem_grant_ready),
    .io_mem_grant_valid(icache_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(icache_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(icache_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(icache_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(icache_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(icache_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(icache_io_mem_grant_bits_data)
  );
  TLB tlb (
    .clk(tlb_clk),
    .reset(tlb_reset),
    .io_req_ready(tlb_io_req_ready),
    .io_req_valid(tlb_io_req_valid),
    .io_req_bits_vpn(tlb_io_req_bits_vpn),
    .io_req_bits_passthrough(tlb_io_req_bits_passthrough),
    .io_req_bits_instruction(tlb_io_req_bits_instruction),
    .io_req_bits_store(tlb_io_req_bits_store),
    .io_resp_miss(tlb_io_resp_miss),
    .io_resp_ppn(tlb_io_resp_ppn),
    .io_resp_xcpt_ld(tlb_io_resp_xcpt_ld),
    .io_resp_xcpt_st(tlb_io_resp_xcpt_st),
    .io_resp_xcpt_if(tlb_io_resp_xcpt_if),
    .io_resp_cacheable(tlb_io_resp_cacheable),
    .io_ptw_req_ready(tlb_io_ptw_req_ready),
    .io_ptw_req_valid(tlb_io_ptw_req_valid),
    .io_ptw_req_bits_prv(tlb_io_ptw_req_bits_prv),
    .io_ptw_req_bits_pum(tlb_io_ptw_req_bits_pum),
    .io_ptw_req_bits_mxr(tlb_io_ptw_req_bits_mxr),
    .io_ptw_req_bits_addr(tlb_io_ptw_req_bits_addr),
    .io_ptw_req_bits_store(tlb_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(tlb_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(tlb_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_reserved_for_hardware(tlb_io_ptw_resp_bits_pte_reserved_for_hardware),
    .io_ptw_resp_bits_pte_ppn(tlb_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(tlb_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(tlb_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(tlb_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(tlb_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(tlb_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(tlb_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(tlb_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(tlb_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(tlb_io_ptw_resp_bits_pte_v),
    .io_ptw_ptbr_asid(tlb_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(tlb_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(tlb_io_ptw_invalidate),
    .io_ptw_status_debug(tlb_io_ptw_status_debug),
    .io_ptw_status_prv(tlb_io_ptw_status_prv),
    .io_ptw_status_sd(tlb_io_ptw_status_sd),
    .io_ptw_status_zero3(tlb_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(tlb_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(tlb_io_ptw_status_zero2),
    .io_ptw_status_vm(tlb_io_ptw_status_vm),
    .io_ptw_status_zero1(tlb_io_ptw_status_zero1),
    .io_ptw_status_mxr(tlb_io_ptw_status_mxr),
    .io_ptw_status_pum(tlb_io_ptw_status_pum),
    .io_ptw_status_mprv(tlb_io_ptw_status_mprv),
    .io_ptw_status_xs(tlb_io_ptw_status_xs),
    .io_ptw_status_fs(tlb_io_ptw_status_fs),
    .io_ptw_status_mpp(tlb_io_ptw_status_mpp),
    .io_ptw_status_hpp(tlb_io_ptw_status_hpp),
    .io_ptw_status_spp(tlb_io_ptw_status_spp),
    .io_ptw_status_mpie(tlb_io_ptw_status_mpie),
    .io_ptw_status_hpie(tlb_io_ptw_status_hpie),
    .io_ptw_status_spie(tlb_io_ptw_status_spie),
    .io_ptw_status_upie(tlb_io_ptw_status_upie),
    .io_ptw_status_mie(tlb_io_ptw_status_mie),
    .io_ptw_status_hie(tlb_io_ptw_status_hie),
    .io_ptw_status_sie(tlb_io_ptw_status_sie),
    .io_ptw_status_uie(tlb_io_ptw_status_uie)
  );
  assign io_cpu_resp_valid = T_1404;
  assign io_cpu_resp_bits_pc = s2_pc;
  assign io_cpu_resp_bits_data_0 = T_1408;
  assign io_cpu_resp_bits_mask = T_1411[0];
  assign io_cpu_resp_bits_xcpt_if = s2_xcpt_if;
  assign io_cpu_resp_bits_replay = T_1417;
  assign io_cpu_btb_resp_valid = s2_btb_resp_valid;
  assign io_cpu_btb_resp_bits_taken = s2_btb_resp_bits_taken;
  assign io_cpu_btb_resp_bits_mask = s2_btb_resp_bits_mask;
  assign io_cpu_btb_resp_bits_bridx = s2_btb_resp_bits_bridx;
  assign io_cpu_btb_resp_bits_target = s2_btb_resp_bits_target;
  assign io_cpu_btb_resp_bits_entry = s2_btb_resp_bits_entry;
  assign io_cpu_btb_resp_bits_bht_history = s2_btb_resp_bits_bht_history;
  assign io_cpu_btb_resp_bits_bht_value = s2_btb_resp_bits_bht_value;
  assign io_cpu_npc = T_1405;
  assign io_ptw_req_valid = tlb_io_ptw_req_valid;
  assign io_ptw_req_bits_prv = tlb_io_ptw_req_bits_prv;
  assign io_ptw_req_bits_pum = tlb_io_ptw_req_bits_pum;
  assign io_ptw_req_bits_mxr = tlb_io_ptw_req_bits_mxr;
  assign io_ptw_req_bits_addr = tlb_io_ptw_req_bits_addr;
  assign io_ptw_req_bits_store = tlb_io_ptw_req_bits_store;
  assign io_ptw_req_bits_fetch = tlb_io_ptw_req_bits_fetch;
  assign io_mem_acquire_valid = icache_io_mem_acquire_valid;
  assign io_mem_acquire_bits_addr_block = icache_io_mem_acquire_bits_addr_block;
  assign io_mem_acquire_bits_client_xact_id = icache_io_mem_acquire_bits_client_xact_id;
  assign io_mem_acquire_bits_addr_beat = icache_io_mem_acquire_bits_addr_beat;
  assign io_mem_acquire_bits_is_builtin_type = icache_io_mem_acquire_bits_is_builtin_type;
  assign io_mem_acquire_bits_a_type = icache_io_mem_acquire_bits_a_type;
  assign io_mem_acquire_bits_union = icache_io_mem_acquire_bits_union;
  assign io_mem_acquire_bits_data = icache_io_mem_acquire_bits_data;
  assign io_mem_grant_ready = icache_io_mem_grant_ready;
  assign icache_clk = clk;
  assign icache_reset = reset;
  assign icache_io_req_valid = T_1392;
  assign icache_io_req_bits_addr = io_cpu_npc;
  assign icache_io_s1_ppn = tlb_io_resp_ppn;
  assign icache_io_s1_kill = T_1396;
  assign icache_io_s2_kill = s2_speculative;
  assign icache_io_resp_ready = T_1401;
  assign icache_io_invalidate = io_cpu_flush_icache;
  assign icache_io_mem_acquire_ready = io_mem_acquire_ready;
  assign icache_io_mem_grant_valid = io_mem_grant_valid;
  assign icache_io_mem_grant_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign icache_io_mem_grant_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign icache_io_mem_grant_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign icache_io_mem_grant_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign icache_io_mem_grant_bits_g_type = io_mem_grant_bits_g_type;
  assign icache_io_mem_grant_bits_data = io_mem_grant_bits_data;
  assign tlb_clk = clk;
  assign tlb_reset = reset;
  assign tlb_io_req_valid = T_1383;
  assign tlb_io_req_bits_vpn = T_1384;
  assign tlb_io_req_bits_passthrough = 1'h0;
  assign tlb_io_req_bits_instruction = 1'h1;
  assign tlb_io_req_bits_store = 1'h0;
  assign tlb_io_ptw_req_ready = io_ptw_req_ready;
  assign tlb_io_ptw_resp_valid = io_ptw_resp_valid;
  assign tlb_io_ptw_resp_bits_pte_reserved_for_hardware = io_ptw_resp_bits_pte_reserved_for_hardware;
  assign tlb_io_ptw_resp_bits_pte_ppn = io_ptw_resp_bits_pte_ppn;
  assign tlb_io_ptw_resp_bits_pte_reserved_for_software = io_ptw_resp_bits_pte_reserved_for_software;
  assign tlb_io_ptw_resp_bits_pte_d = io_ptw_resp_bits_pte_d;
  assign tlb_io_ptw_resp_bits_pte_a = io_ptw_resp_bits_pte_a;
  assign tlb_io_ptw_resp_bits_pte_g = io_ptw_resp_bits_pte_g;
  assign tlb_io_ptw_resp_bits_pte_u = io_ptw_resp_bits_pte_u;
  assign tlb_io_ptw_resp_bits_pte_x = io_ptw_resp_bits_pte_x;
  assign tlb_io_ptw_resp_bits_pte_w = io_ptw_resp_bits_pte_w;
  assign tlb_io_ptw_resp_bits_pte_r = io_ptw_resp_bits_pte_r;
  assign tlb_io_ptw_resp_bits_pte_v = io_ptw_resp_bits_pte_v;
  assign tlb_io_ptw_ptbr_asid = io_ptw_ptbr_asid;
  assign tlb_io_ptw_ptbr_ppn = io_ptw_ptbr_ppn;
  assign tlb_io_ptw_invalidate = io_ptw_invalidate;
  assign tlb_io_ptw_status_debug = io_ptw_status_debug;
  assign tlb_io_ptw_status_prv = io_ptw_status_prv;
  assign tlb_io_ptw_status_sd = io_ptw_status_sd;
  assign tlb_io_ptw_status_zero3 = io_ptw_status_zero3;
  assign tlb_io_ptw_status_sd_rv32 = io_ptw_status_sd_rv32;
  assign tlb_io_ptw_status_zero2 = io_ptw_status_zero2;
  assign tlb_io_ptw_status_vm = io_ptw_status_vm;
  assign tlb_io_ptw_status_zero1 = io_ptw_status_zero1;
  assign tlb_io_ptw_status_mxr = io_ptw_status_mxr;
  assign tlb_io_ptw_status_pum = io_ptw_status_pum;
  assign tlb_io_ptw_status_mprv = io_ptw_status_mprv;
  assign tlb_io_ptw_status_xs = io_ptw_status_xs;
  assign tlb_io_ptw_status_fs = io_ptw_status_fs;
  assign tlb_io_ptw_status_mpp = io_ptw_status_mpp;
  assign tlb_io_ptw_status_hpp = io_ptw_status_hpp;
  assign tlb_io_ptw_status_spp = io_ptw_status_spp;
  assign tlb_io_ptw_status_mpie = io_ptw_status_mpie;
  assign tlb_io_ptw_status_hpie = io_ptw_status_hpie;
  assign tlb_io_ptw_status_spie = io_ptw_status_spie;
  assign tlb_io_ptw_status_upie = io_ptw_status_upie;
  assign tlb_io_ptw_status_mie = io_ptw_status_mie;
  assign tlb_io_ptw_status_hie = io_ptw_status_hie;
  assign tlb_io_ptw_status_sie = io_ptw_status_sie;
  assign tlb_io_ptw_status_uie = io_ptw_status_uie;
  assign T_1315 = ~ s1_pc_;
  assign T_1317 = T_1315 | 32'h3;
  assign s1_pc = ~ T_1317;
  assign T_1342 = ~ s1_pc;
  assign T_1344 = T_1342 | 32'h3;
  assign T_1345 = ~ T_1344;
  assign T_1347 = T_1345 + 32'h4;
  assign ntpc = T_1347[31:0];
  assign predicted_npc = ntpc;
  assign T_1349 = icache_io_resp_valid == 1'h0;
  assign icmiss = s2_valid & T_1349;
  assign npc = icmiss ? s2_pc : predicted_npc;
  assign T_1351 = icmiss == 1'h0;
  assign T_1353 = io_cpu_req_valid == 1'h0;
  assign T_1354 = T_1351 & T_1353;
  assign T_1356 = ntpc & 32'h8;
  assign T_1358 = s1_pc & 32'h8;
  assign T_1359 = T_1356 == T_1358;
  assign T_1360 = T_1354 & T_1359;
  assign s0_same_block = T_1360;
  assign T_1362 = io_cpu_resp_ready == 1'h0;
  assign stall = io_cpu_resp_valid & T_1362;
  assign T_1364 = stall == 1'h0;
  assign T_1366 = tlb_io_resp_miss == 1'h0;
  assign T_1367 = s0_same_block & T_1366;
  assign T_1369 = icmiss ? s2_speculative : 1'h1;
  assign T_1375 = tlb_io_resp_cacheable == 1'h0;
  assign T_1376 = s1_speculative & T_1375;
  assign GEN_0 = T_1351 ? s1_pc : s2_pc;
  assign GEN_1 = T_1351 ? T_1376 : s2_speculative;
  assign GEN_2 = T_1351 ? tlb_io_resp_xcpt_if : s2_xcpt_if;
  assign GEN_3 = T_1364 ? T_1367 : s1_same_block;
  assign GEN_4 = T_1364 ? npc : s1_pc_;
  assign GEN_5 = T_1364 ? T_1369 : s1_speculative;
  assign GEN_6 = T_1364 ? T_1351 : s2_valid;
  assign GEN_7 = T_1364 ? GEN_0 : s2_pc;
  assign GEN_8 = T_1364 ? GEN_1 : s2_speculative;
  assign GEN_9 = T_1364 ? GEN_2 : s2_xcpt_if;
  assign GEN_10 = io_cpu_req_valid ? 1'h0 : GEN_3;
  assign GEN_11 = io_cpu_req_valid ? io_cpu_req_bits_pc : GEN_4;
  assign GEN_12 = io_cpu_req_valid ? io_cpu_req_bits_speculative : GEN_5;
  assign GEN_13 = io_cpu_req_valid ? 1'h0 : GEN_6;
  assign T_1383 = T_1364 & T_1351;
  assign T_1384 = s1_pc[31:12];
  assign T_1391 = s0_same_block == 1'h0;
  assign T_1392 = T_1364 & T_1391;
  assign T_1393 = io_cpu_req_valid | tlb_io_resp_miss;
  assign T_1394 = T_1393 | tlb_io_resp_xcpt_if;
  assign T_1395 = T_1394 | icmiss;
  assign T_1396 = T_1395 | io_cpu_flush_tlb;
  assign T_1400 = s1_same_block == 1'h0;
  assign T_1401 = T_1364 & T_1400;
  assign T_1402 = icache_io_resp_valid | s2_speculative;
  assign T_1403 = T_1402 | s2_xcpt_if;
  assign T_1404 = s2_valid & T_1403;
  assign T_1405 = io_cpu_req_valid ? io_cpu_req_bits_pc : npc;
  assign T_1406 = s2_pc[2];
  assign GEN_14 = {{5'd0}, T_1406};
  assign T_1407 = GEN_14 << 5;
  assign fetch_data = icache_io_resp_bits_datablock >> T_1407;
  assign T_1408 = fetch_data[31:0];
  assign T_1411 = 2'h1 << T_1406;
  assign T_1414 = s2_speculative & T_1349;
  assign T_1416 = s2_xcpt_if == 1'h0;
  assign T_1417 = T_1414 & T_1416;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_15 = {1{$random}};
  s1_pc_ = GEN_15[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_16 = {1{$random}};
  s1_speculative = GEN_16[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_17 = {1{$random}};
  s1_same_block = GEN_17[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_18 = {1{$random}};
  s2_valid = GEN_18[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_19 = {1{$random}};
  s2_pc = GEN_19[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_20 = {1{$random}};
  s2_btb_resp_valid = GEN_20[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_21 = {1{$random}};
  s2_btb_resp_bits_taken = GEN_21[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_22 = {1{$random}};
  s2_btb_resp_bits_mask = GEN_22[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_23 = {1{$random}};
  s2_btb_resp_bits_bridx = GEN_23[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_24 = {1{$random}};
  s2_btb_resp_bits_target = GEN_24[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_25 = {1{$random}};
  s2_btb_resp_bits_entry = GEN_25[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_26 = {1{$random}};
  s2_btb_resp_bits_bht_history = GEN_26[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_27 = {1{$random}};
  s2_btb_resp_bits_bht_value = GEN_27[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_28 = {1{$random}};
  s2_xcpt_if = GEN_28[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_29 = {1{$random}};
  s2_speculative = GEN_29[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(io_cpu_req_valid) begin
        s1_pc_ <= io_cpu_req_bits_pc;
      end else begin
        if(T_1364) begin
          if(icmiss) begin
            s1_pc_ <= s2_pc;
          end else begin
            s1_pc_ <= predicted_npc;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_cpu_req_valid) begin
        s1_speculative <= io_cpu_req_bits_speculative;
      end else begin
        if(T_1364) begin
          if(icmiss) begin
            s1_speculative <= s2_speculative;
          end else begin
            s1_speculative <= 1'h1;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(io_cpu_req_valid) begin
        s1_same_block <= 1'h0;
      end else begin
        if(T_1364) begin
          s1_same_block <= T_1367;
        end
      end
    end
    if(reset) begin
      s2_valid <= 1'h1;
    end else begin
      if(io_cpu_req_valid) begin
        s2_valid <= 1'h0;
      end else begin
        if(T_1364) begin
          s2_valid <= T_1351;
        end
      end
    end
    if(reset) begin
//<CJ>      s2_pc <= 32'h60000000;
      s2_pc <= RESET_VECTOR_ADDR;
    end else begin
      if(T_1364) begin
        if(T_1351) begin
          s2_pc <= s1_pc;
        end
      end
    end
    if(reset) begin
      s2_btb_resp_valid <= 1'h0;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(reset) begin
      s2_xcpt_if <= 1'h0;
    end else begin
      if(T_1364) begin
        if(T_1351) begin
          s2_xcpt_if <= tlb_io_resp_xcpt_if;
        end
      end
    end
    if(reset) begin
      s2_speculative <= 1'h0;
    end else begin
      if(T_1364) begin
        if(T_1351) begin
          s2_speculative <= T_1376;
        end
      end
    end
  end
endmodule
module FinishQueue(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_manager_xact_id,
  input   io_enq_bits_manager_id,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_manager_xact_id,
  output  io_deq_bits_manager_id,
  output  io_count
);
  reg [1:0] ram_manager_xact_id [0:0];
  reg [31:0] GEN_0;
  wire [1:0] ram_manager_xact_id_T_254_data;
  wire  ram_manager_xact_id_T_254_addr;
  wire  ram_manager_xact_id_T_254_en;
  wire [1:0] ram_manager_xact_id_T_224_data;
  wire  ram_manager_xact_id_T_224_addr;
  wire  ram_manager_xact_id_T_224_mask;
  wire  ram_manager_xact_id_T_224_en;
  reg  ram_manager_id [0:0];
  reg [31:0] GEN_1;
  wire  ram_manager_id_T_254_data;
  wire  ram_manager_id_T_254_addr;
  wire  ram_manager_id_T_254_en;
  wire  ram_manager_id_T_224_data;
  wire  ram_manager_id_T_224_addr;
  wire  ram_manager_id_T_224_mask;
  wire  ram_manager_id_T_224_en;
  reg  maybe_full;
  reg [31:0] GEN_2;
  wire  T_221;
  wire  T_222;
  wire  do_enq;
  wire  T_223;
  wire  do_deq;
  wire  T_249;
  wire  GEN_7;
  wire  T_251;
  wire [1:0] T_277;
  wire  ptr_diff;
  wire [1:0] T_279;
  assign io_enq_ready = T_221;
  assign io_deq_valid = T_251;
  assign io_deq_bits_manager_xact_id = ram_manager_xact_id_T_254_data;
  assign io_deq_bits_manager_id = ram_manager_id_T_254_data;
  assign io_count = T_279[0];
  assign ram_manager_xact_id_T_254_addr = 1'h0;
  assign ram_manager_xact_id_T_254_en = 1'h1;
  assign ram_manager_xact_id_T_254_data = ram_manager_xact_id[ram_manager_xact_id_T_254_addr];
  assign ram_manager_xact_id_T_224_data = io_enq_bits_manager_xact_id;
  assign ram_manager_xact_id_T_224_addr = 1'h0;
  assign ram_manager_xact_id_T_224_mask = do_enq;
  assign ram_manager_xact_id_T_224_en = do_enq;
  assign ram_manager_id_T_254_addr = 1'h0;
  assign ram_manager_id_T_254_en = 1'h1;
  assign ram_manager_id_T_254_data = ram_manager_id[ram_manager_id_T_254_addr];
  assign ram_manager_id_T_224_data = io_enq_bits_manager_id;
  assign ram_manager_id_T_224_addr = 1'h0;
  assign ram_manager_id_T_224_mask = do_enq;
  assign ram_manager_id_T_224_en = do_enq;
  assign T_221 = maybe_full == 1'h0;
  assign T_222 = io_enq_ready & io_enq_valid;
  assign do_enq = T_222;
  assign T_223 = io_deq_ready & io_deq_valid;
  assign do_deq = T_223;
  assign T_249 = do_enq != do_deq;
  assign GEN_7 = T_249 ? do_enq : maybe_full;
  assign T_251 = T_221 == 1'h0;
  assign T_277 = 1'h0 - 1'h0;
  assign ptr_diff = T_277[0:0];
  assign T_279 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_manager_xact_id[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_manager_id[initvar] = GEN_1[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_2 = {1{$random}};
  maybe_full = GEN_2[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_manager_xact_id_T_224_en & ram_manager_xact_id_T_224_mask) begin
      ram_manager_xact_id[ram_manager_xact_id_T_224_addr] <= ram_manager_xact_id_T_224_data;
    end
    if(ram_manager_id_T_224_en & ram_manager_id_T_224_mask) begin
      ram_manager_id[ram_manager_id_T_224_addr] <= ram_manager_id_T_224_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_249) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module MetadataArray(
  input   clk,
  input   reset,
  output  io_read_ready,
  input   io_read_valid,
  input  [6:0] io_read_bits_idx,
  input   io_read_bits_way_en,
  output  io_write_ready,
  input   io_write_valid,
  input  [6:0] io_write_bits_idx,
  input   io_write_bits_way_en,
  input  [18:0] io_write_bits_data_tag,
  input  [1:0] io_write_bits_data_coh_state,
  output [18:0] io_resp_0_tag,
  output [1:0] io_resp_0_coh_state
);
  wire [1:0] T_44_state;
  wire [18:0] rstVal_tag;
  wire [1:0] rstVal_coh_state;
  reg [7:0] rst_cnt;
  reg [31:0] GEN_1;
  wire  rst;
  wire [7:0] waddr;
  wire [18:0] T_1569_tag;
  wire [1:0] T_1569_coh_state;
  wire [20:0] wdata;
  wire [8:0] T_1666;
  wire [7:0] T_1667;
  wire [7:0] GEN_0;
  reg [20:0] T_1676_0 [0:127];
  reg [31:0] GEN_2;
  wire [20:0] T_1676_0_T_1693_data;
  wire [6:0] T_1676_0_T_1693_addr;
  wire  T_1676_0_T_1693_en;
  reg [6:0] GEN_3;
  reg [31:0] GEN_4;
  reg  GEN_5;
  reg [31:0] GEN_6;
  wire [20:0] T_1676_0_T_1687_data;
  wire [6:0] T_1676_0_T_1687_addr;
  wire  T_1676_0_T_1687_mask;
  wire  T_1676_0_T_1687_en;
  wire  T_1677;
  wire [20:0] T_1683_0;
  wire [6:0] T_1690;
  wire [18:0] T_2199_0_tag;
  wire [1:0] T_2199_0_coh_state;
  wire [1:0] T_2367;
  wire [18:0] T_2368;
  wire  T_2370;
  wire  T_2372;
  wire  T_2373;
  assign io_read_ready = T_2373;
  assign io_write_ready = T_2370;
  assign io_resp_0_tag = T_2199_0_tag;
  assign io_resp_0_coh_state = T_2199_0_coh_state;
  assign T_44_state = 2'h0;
  assign rstVal_tag = 19'h0;
  assign rstVal_coh_state = T_44_state;
  assign rst = rst_cnt < 8'h80;
  assign waddr = rst ? rst_cnt : {{1'd0}, io_write_bits_idx};
  assign T_1569_tag = rst ? rstVal_tag : io_write_bits_data_tag;
  assign T_1569_coh_state = rst ? rstVal_coh_state : io_write_bits_data_coh_state;
  assign wdata = {T_1569_tag,T_1569_coh_state};
  assign T_1666 = rst_cnt + 8'h1;
  assign T_1667 = T_1666[7:0];
  assign GEN_0 = rst ? T_1667 : rst_cnt;
  assign T_1676_0_T_1693_addr = T_1690;
  assign T_1676_0_T_1693_en = 1'h1;
  assign T_1676_0_T_1693_data = T_1676_0[GEN_3];
  assign T_1676_0_T_1687_data = T_1683_0;
  assign T_1676_0_T_1687_addr = waddr[6:0];
  assign T_1676_0_T_1687_mask = T_1677;
  assign T_1676_0_T_1687_en = T_1677;
  assign T_1677 = rst | io_write_valid;
  assign T_1683_0 = wdata;
  assign T_1690 = io_read_bits_idx;
  assign T_2199_0_tag = T_2368;
  assign T_2199_0_coh_state = T_2367;
  assign T_2367 = T_1676_0_T_1693_data[1:0];
  assign T_2368 = T_1676_0_T_1693_data[20:2];
  assign T_2370 = rst == 1'h0;
  assign T_2372 = io_write_valid == 1'h0;
  assign T_2373 = T_2370 & T_2372;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_1 = {1{$random}};
  rst_cnt = GEN_1[7:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    T_1676_0[initvar] = GEN_2[20:0];
  `endif
  `ifdef RANDOMIZE
  GEN_4 = {1{$random}};
  GEN_3 = GEN_4[6:0];
  `endif
  `ifdef RANDOMIZE
  GEN_6 = {1{$random}};
  GEN_5 = GEN_6[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      rst_cnt <= 8'h0;
    end else begin
      if(rst) begin
        rst_cnt <= T_1667;
      end
    end
    GEN_3 <= T_1676_0_T_1693_addr;
    GEN_5 <= T_1676_0_T_1693_en;
    if(T_1676_0_T_1687_en & T_1676_0_T_1687_mask) begin
      T_1676_0[T_1676_0_T_1687_addr] <= T_1676_0_T_1687_data;
    end
  end
endmodule
module Arbiter(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [6:0] io_in_0_bits_idx,
  input   io_in_0_bits_way_en,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [6:0] io_in_1_bits_idx,
  input   io_in_1_bits_way_en,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [6:0] io_in_2_bits_idx,
  input   io_in_2_bits_way_en,
  input   io_out_ready,
  output  io_out_valid,
  output [6:0] io_out_bits_idx,
  output  io_out_bits_way_en,
  output [1:0] io_chosen
);
  wire [1:0] GEN_0;
  wire [6:0] GEN_1;
  wire  GEN_2;
  wire [1:0] GEN_3;
  wire [6:0] GEN_4;
  wire  GEN_5;
  wire  T_638;
  wire  T_640;
  wire  T_642;
  wire  T_644;
  wire  T_645;
  wire  T_647;
  wire  T_648;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_644;
  assign io_in_2_ready = T_645;
  assign io_out_valid = T_648;
  assign io_out_bits_idx = GEN_4;
  assign io_out_bits_way_en = GEN_5;
  assign io_chosen = GEN_3;
  assign GEN_0 = io_in_1_valid ? 2'h1 : 2'h2;
  assign GEN_1 = io_in_1_valid ? io_in_1_bits_idx : io_in_2_bits_idx;
  assign GEN_2 = io_in_1_valid ? io_in_1_bits_way_en : io_in_2_bits_way_en;
  assign GEN_3 = io_in_0_valid ? 2'h0 : GEN_0;
  assign GEN_4 = io_in_0_valid ? io_in_0_bits_idx : GEN_1;
  assign GEN_5 = io_in_0_valid ? io_in_0_bits_way_en : GEN_2;
  assign T_638 = io_in_0_valid | io_in_1_valid;
  assign T_640 = io_in_0_valid == 1'h0;
  assign T_642 = T_638 == 1'h0;
  assign T_644 = T_640 & io_out_ready;
  assign T_645 = T_642 & io_out_ready;
  assign T_647 = T_642 == 1'h0;
  assign T_648 = T_647 | io_in_2_valid;
endmodule
module Arbiter_1(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [6:0] io_in_0_bits_idx,
  input   io_in_0_bits_way_en,
  input  [18:0] io_in_0_bits_data_tag,
  input  [1:0] io_in_0_bits_data_coh_state,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [6:0] io_in_1_bits_idx,
  input   io_in_1_bits_way_en,
  input  [18:0] io_in_1_bits_data_tag,
  input  [1:0] io_in_1_bits_data_coh_state,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [6:0] io_in_2_bits_idx,
  input   io_in_2_bits_way_en,
  input  [18:0] io_in_2_bits_data_tag,
  input  [1:0] io_in_2_bits_data_coh_state,
  input   io_out_ready,
  output  io_out_valid,
  output [6:0] io_out_bits_idx,
  output  io_out_bits_way_en,
  output [18:0] io_out_bits_data_tag,
  output [1:0] io_out_bits_data_coh_state,
  output [1:0] io_chosen
);
  wire [1:0] GEN_0;
  wire [6:0] GEN_1;
  wire  GEN_2;
  wire [18:0] GEN_3;
  wire [1:0] GEN_4;
  wire [1:0] GEN_5;
  wire [6:0] GEN_6;
  wire  GEN_7;
  wire [18:0] GEN_8;
  wire [1:0] GEN_9;
  wire  T_2822;
  wire  T_2824;
  wire  T_2826;
  wire  T_2828;
  wire  T_2829;
  wire  T_2831;
  wire  T_2832;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_2828;
  assign io_in_2_ready = T_2829;
  assign io_out_valid = T_2832;
  assign io_out_bits_idx = GEN_6;
  assign io_out_bits_way_en = GEN_7;
  assign io_out_bits_data_tag = GEN_8;
  assign io_out_bits_data_coh_state = GEN_9;
  assign io_chosen = GEN_5;
  assign GEN_0 = io_in_1_valid ? 2'h1 : 2'h2;
  assign GEN_1 = io_in_1_valid ? io_in_1_bits_idx : io_in_2_bits_idx;
  assign GEN_2 = io_in_1_valid ? io_in_1_bits_way_en : io_in_2_bits_way_en;
  assign GEN_3 = io_in_1_valid ? io_in_1_bits_data_tag : io_in_2_bits_data_tag;
  assign GEN_4 = io_in_1_valid ? io_in_1_bits_data_coh_state : io_in_2_bits_data_coh_state;
  assign GEN_5 = io_in_0_valid ? 2'h0 : GEN_0;
  assign GEN_6 = io_in_0_valid ? io_in_0_bits_idx : GEN_1;
  assign GEN_7 = io_in_0_valid ? io_in_0_bits_way_en : GEN_2;
  assign GEN_8 = io_in_0_valid ? io_in_0_bits_data_tag : GEN_3;
  assign GEN_9 = io_in_0_valid ? io_in_0_bits_data_coh_state : GEN_4;
  assign T_2822 = io_in_0_valid | io_in_1_valid;
  assign T_2824 = io_in_0_valid == 1'h0;
  assign T_2826 = T_2822 == 1'h0;
  assign T_2828 = T_2824 & io_out_ready;
  assign T_2829 = T_2826 & io_out_ready;
  assign T_2831 = T_2826 == 1'h0;
  assign T_2832 = T_2831 | io_in_2_valid;
endmodule
module DCacheDataArray(
  input   clk,
  input   reset,
  input   io_req_valid,
  input  [12:0] io_req_bits_addr,
  input   io_req_bits_write,
  input  [63:0] io_req_bits_wdata,
  input  [7:0] io_req_bits_wmask,
  input   io_req_bits_way_en,
  output [63:0] io_resp_0
);
  wire [9:0] addr;
  reg [7:0] T_406_0 [0:1023];
  reg [31:0] GEN_0;
  wire [7:0] T_406_0_T_446_data;
  wire [9:0] T_406_0_T_446_addr;
  wire  T_406_0_T_446_en;
  reg [9:0] GEN_1/* synthesis syn_keep=1 */;
  reg [31:0] GEN_2;
  reg  GEN_3;
  reg [31:0] GEN_4;
  wire [7:0] T_406_0_T_437_data;
  wire [9:0] T_406_0_T_437_addr;
  wire  T_406_0_T_437_mask;
  wire  T_406_0_T_437_en;
  reg [7:0] T_406_1 [0:1023];
  reg [31:0] GEN_5;
  wire [7:0] T_406_1_T_446_data;
  wire [9:0] T_406_1_T_446_addr;
  wire  T_406_1_T_446_en;
  reg [9:0] GEN_6/* synthesis syn_keep=1 */;
  reg [31:0] GEN_7;
  reg  GEN_8;
  reg [31:0] GEN_9;
  wire [7:0] T_406_1_T_437_data;
  wire [9:0] T_406_1_T_437_addr;
  wire  T_406_1_T_437_mask;
  wire  T_406_1_T_437_en;
  reg [7:0] T_406_2 [0:1023];
  reg [31:0] GEN_10;
  wire [7:0] T_406_2_T_446_data;
  wire [9:0] T_406_2_T_446_addr;
  wire  T_406_2_T_446_en;
  reg [9:0] GEN_11/* synthesis syn_keep=1 */;
  reg [31:0] GEN_12;
  reg  GEN_13;
  reg [31:0] GEN_14;
  wire [7:0] T_406_2_T_437_data;
  wire [9:0] T_406_2_T_437_addr;
  wire  T_406_2_T_437_mask;
  wire  T_406_2_T_437_en;
  reg [7:0] T_406_3 [0:1023];
  reg [31:0] GEN_15;
  wire [7:0] T_406_3_T_446_data;
  wire [9:0] T_406_3_T_446_addr;
  wire  T_406_3_T_446_en;
  reg [9:0] GEN_16/* synthesis syn_keep=1 */;
  reg [31:0] GEN_17;
  reg  GEN_18;
  reg [31:0] GEN_19;
  wire [7:0] T_406_3_T_437_data;
  wire [9:0] T_406_3_T_437_addr;
  wire  T_406_3_T_437_mask;
  wire  T_406_3_T_437_en;
  reg [7:0] T_406_4 [0:1023];
  reg [31:0] GEN_20;
  wire [7:0] T_406_4_T_446_data;
  wire [9:0] T_406_4_T_446_addr;
  wire  T_406_4_T_446_en;
  reg [9:0] GEN_21/* synthesis syn_keep=1 */;
  reg [31:0] GEN_22;
  reg  GEN_23;
  reg [31:0] GEN_24;
  wire [7:0] T_406_4_T_437_data;
  wire [9:0] T_406_4_T_437_addr;
  wire  T_406_4_T_437_mask;
  wire  T_406_4_T_437_en;
  reg [7:0] T_406_5 [0:1023];
  reg [31:0] GEN_25;
  wire [7:0] T_406_5_T_446_data;
  wire [9:0] T_406_5_T_446_addr;
  wire  T_406_5_T_446_en;
  reg [9:0] GEN_26/* synthesis syn_keep=1 */;
  reg [31:0] GEN_27;
  reg  GEN_29;
  reg [31:0] GEN_31;
  wire [7:0] T_406_5_T_437_data;
  wire [9:0] T_406_5_T_437_addr;
  wire  T_406_5_T_437_mask;
  wire  T_406_5_T_437_en;
  reg [7:0] T_406_6 [0:1023];
  reg [31:0] GEN_33;
  wire [7:0] T_406_6_T_446_data;
  wire [9:0] T_406_6_T_446_addr;
  wire  T_406_6_T_446_en;
  reg [9:0] GEN_35/* synthesis syn_keep=1 */;
  reg [31:0] GEN_37;
  reg  GEN_39;
  reg [31:0] GEN_41;
  wire [7:0] T_406_6_T_437_data;
  wire [9:0] T_406_6_T_437_addr;
  wire  T_406_6_T_437_mask;
  wire  T_406_6_T_437_en;
  reg [7:0] T_406_7 [0:1023];
  reg [31:0] GEN_43;
  wire [7:0] T_406_7_T_446_data;
  wire [9:0] T_406_7_T_446_addr;
  wire  T_406_7_T_446_en;
  reg [9:0] GEN_44/* synthesis syn_keep=1 */;
  reg [31:0] GEN_45;
  reg  GEN_46;
  reg [31:0] GEN_47;
  wire [7:0] T_406_7_T_437_data;
  wire [9:0] T_406_7_T_437_addr;
  wire  T_406_7_T_437_mask;
  wire  T_406_7_T_437_en;
  wire  T_411;
  wire [7:0] T_412;
  wire [7:0] T_413;
  wire [7:0] T_414;
  wire [7:0] T_415;
  wire [7:0] T_416;
  wire [7:0] T_417;
  wire [7:0] T_418;
  wire [7:0] T_419;
  wire [7:0] T_425_0;
  wire [7:0] T_425_1;
  wire [7:0] T_425_2;
  wire [7:0] T_425_3;
  wire [7:0] T_425_4;
  wire [7:0] T_425_5;
  wire [7:0] T_425_6;
  wire [7:0] T_425_7;
  wire  T_427;
  wire  T_428;
  wire  T_429;
  wire  T_430;
  wire  T_431;
  wire  T_432;
  wire  T_433;
  wire  T_434;
  wire  GEN_28;
  wire  GEN_30;
  wire  GEN_32;
  wire  GEN_34;
  wire  GEN_36;
  wire  GEN_38;
  wire  GEN_40;
  wire  GEN_42;
  wire [9:0] T_443;
  wire [15:0] T_448;
  wire [15:0] T_449;
  wire [31:0] T_450;
  wire [15:0] T_451;
  wire [15:0] T_452;
  wire [31:0] T_453;
  wire [63:0] T_454;
  assign io_resp_0 = T_454;
  assign addr = io_req_bits_addr[12:3];
  assign T_406_0_T_446_addr = T_443;
  assign T_406_0_T_446_en = 1'h1;
  assign T_406_0_T_446_data = T_406_0[GEN_1];
  assign T_406_0_T_437_data = T_425_0;
  assign T_406_0_T_437_addr = addr;
  assign T_406_0_T_437_mask = GEN_28;
  assign T_406_0_T_437_en = T_411;
  assign T_406_1_T_446_addr = T_443;
  assign T_406_1_T_446_en = 1'h1;
  assign T_406_1_T_446_data = T_406_1[GEN_6];
  assign T_406_1_T_437_data = T_425_1;
  assign T_406_1_T_437_addr = addr;
  assign T_406_1_T_437_mask = GEN_30;
  assign T_406_1_T_437_en = T_411;
  assign T_406_2_T_446_addr = T_443;
  assign T_406_2_T_446_en = 1'h1;
  assign T_406_2_T_446_data = T_406_2[GEN_11];
  assign T_406_2_T_437_data = T_425_2;
  assign T_406_2_T_437_addr = addr;
  assign T_406_2_T_437_mask = GEN_32;
  assign T_406_2_T_437_en = T_411;
  assign T_406_3_T_446_addr = T_443;
  assign T_406_3_T_446_en = 1'h1;
  assign T_406_3_T_446_data = T_406_3[GEN_16];
  assign T_406_3_T_437_data = T_425_3;
  assign T_406_3_T_437_addr = addr;
  assign T_406_3_T_437_mask = GEN_34;
  assign T_406_3_T_437_en = T_411;
  assign T_406_4_T_446_addr = T_443;
  assign T_406_4_T_446_en = 1'h1;
  assign T_406_4_T_446_data = T_406_4[GEN_21];
  assign T_406_4_T_437_data = T_425_4;
  assign T_406_4_T_437_addr = addr;
  assign T_406_4_T_437_mask = GEN_36;
  assign T_406_4_T_437_en = T_411;
  assign T_406_5_T_446_addr = T_443;
  assign T_406_5_T_446_en = 1'h1;
  assign T_406_5_T_446_data = T_406_5[GEN_26];
  assign T_406_5_T_437_data = T_425_5;
  assign T_406_5_T_437_addr = addr;
  assign T_406_5_T_437_mask = GEN_38;
  assign T_406_5_T_437_en = T_411;
  assign T_406_6_T_446_addr = T_443;
  assign T_406_6_T_446_en = 1'h1;
  assign T_406_6_T_446_data = T_406_6[GEN_35];
  assign T_406_6_T_437_data = T_425_6;
  assign T_406_6_T_437_addr = addr;
  assign T_406_6_T_437_mask = GEN_40;
  assign T_406_6_T_437_en = T_411;
  assign T_406_7_T_446_addr = T_443;
  assign T_406_7_T_446_en = 1'h1;
  assign T_406_7_T_446_data = T_406_7[GEN_44];
  assign T_406_7_T_437_data = T_425_7;
  assign T_406_7_T_437_addr = addr;
  assign T_406_7_T_437_mask = GEN_42;
  assign T_406_7_T_437_en = T_411;
  assign T_411 = io_req_valid & io_req_bits_write;
  assign T_412 = io_req_bits_wdata[7:0];
  assign T_413 = io_req_bits_wdata[15:8];
  assign T_414 = io_req_bits_wdata[23:16];
  assign T_415 = io_req_bits_wdata[31:24];
  assign T_416 = io_req_bits_wdata[39:32];
  assign T_417 = io_req_bits_wdata[47:40];
  assign T_418 = io_req_bits_wdata[55:48];
  assign T_419 = io_req_bits_wdata[63:56];
  assign T_425_0 = T_412;
  assign T_425_1 = T_413;
  assign T_425_2 = T_414;
  assign T_425_3 = T_415;
  assign T_425_4 = T_416;
  assign T_425_5 = T_417;
  assign T_425_6 = T_418;
  assign T_425_7 = T_419;
  assign T_427 = io_req_bits_wmask[0];
  assign T_428 = io_req_bits_wmask[1];
  assign T_429 = io_req_bits_wmask[2];
  assign T_430 = io_req_bits_wmask[3];
  assign T_431 = io_req_bits_wmask[4];
  assign T_432 = io_req_bits_wmask[5];
  assign T_433 = io_req_bits_wmask[6];
  assign T_434 = io_req_bits_wmask[7];
  assign GEN_28 = T_411 ? T_427 : 1'h0;
  assign GEN_30 = T_411 ? T_428 : 1'h0;
  assign GEN_32 = T_411 ? T_429 : 1'h0;
  assign GEN_34 = T_411 ? T_430 : 1'h0;
  assign GEN_36 = T_411 ? T_431 : 1'h0;
  assign GEN_38 = T_411 ? T_432 : 1'h0;
  assign GEN_40 = T_411 ? T_433 : 1'h0;
  assign GEN_42 = T_411 ? T_434 : 1'h0;
  assign T_443 = addr;
  assign T_448 = {T_406_1_T_446_data,T_406_0_T_446_data};
  assign T_449 = {T_406_3_T_446_data,T_406_2_T_446_data};
  assign T_450 = {T_449,T_448};
  assign T_451 = {T_406_5_T_446_data,T_406_4_T_446_data};
  assign T_452 = {T_406_7_T_446_data,T_406_6_T_446_data};
  assign T_453 = {T_452,T_451};
  assign T_454 = {T_453,T_450};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    T_406_0[initvar] = GEN_0[7:0];
  `endif
  `ifdef RANDOMIZE
  GEN_2 = {1{$random}};
  GEN_1 = GEN_2[9:0];
  `endif
  `ifdef RANDOMIZE
  GEN_4 = {1{$random}};
  GEN_3 = GEN_4[0:0];
  `endif
  GEN_5 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    T_406_1[initvar] = GEN_5[7:0];
  `endif
  `ifdef RANDOMIZE
  GEN_7 = {1{$random}};
  GEN_6 = GEN_7[9:0];
  `endif
  `ifdef RANDOMIZE
  GEN_9 = {1{$random}};
  GEN_8 = GEN_9[0:0];
  `endif
  GEN_10 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    T_406_2[initvar] = GEN_10[7:0];
  `endif
  `ifdef RANDOMIZE
  GEN_12 = {1{$random}};
  GEN_11 = GEN_12[9:0];
  `endif
  `ifdef RANDOMIZE
  GEN_14 = {1{$random}};
  GEN_13 = GEN_14[0:0];
  `endif
  GEN_15 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    T_406_3[initvar] = GEN_15[7:0];
  `endif
  `ifdef RANDOMIZE
  GEN_17 = {1{$random}};
  GEN_16 = GEN_17[9:0];
  `endif
  `ifdef RANDOMIZE
  GEN_19 = {1{$random}};
  GEN_18 = GEN_19[0:0];
  `endif
  GEN_20 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    T_406_4[initvar] = GEN_20[7:0];
  `endif
  `ifdef RANDOMIZE
  GEN_22 = {1{$random}};
  GEN_21 = GEN_22[9:0];
  `endif
  `ifdef RANDOMIZE
  GEN_24 = {1{$random}};
  GEN_23 = GEN_24[0:0];
  `endif
  GEN_25 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    T_406_5[initvar] = GEN_25[7:0];
  `endif
  `ifdef RANDOMIZE
  GEN_27 = {1{$random}};
  GEN_26 = GEN_27[9:0];
  `endif
  `ifdef RANDOMIZE
  GEN_31 = {1{$random}};
  GEN_29 = GEN_31[0:0];
  `endif
  GEN_33 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    T_406_6[initvar] = GEN_33[7:0];
  `endif
  `ifdef RANDOMIZE
  GEN_37 = {1{$random}};
  GEN_35 = GEN_37[9:0];
  `endif
  `ifdef RANDOMIZE
  GEN_41 = {1{$random}};
  GEN_39 = GEN_41[0:0];
  `endif
  GEN_43 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    T_406_7[initvar] = GEN_43[7:0];
  `endif
  `ifdef RANDOMIZE
  GEN_45 = {1{$random}};
  GEN_44 = GEN_45[9:0];
  `endif
  `ifdef RANDOMIZE
  GEN_47 = {1{$random}};
  GEN_46 = GEN_47[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    GEN_1 <= T_406_0_T_446_addr;
    GEN_3 <= T_406_0_T_446_en;
    if(T_406_0_T_437_en & T_406_0_T_437_mask) begin
      T_406_0[T_406_0_T_437_addr] <= T_406_0_T_437_data;
    end
    GEN_6 <= T_406_1_T_446_addr;
    GEN_8 <= T_406_1_T_446_en;
    if(T_406_1_T_437_en & T_406_1_T_437_mask) begin
      T_406_1[T_406_1_T_437_addr] <= T_406_1_T_437_data;
    end
    GEN_11 <= T_406_2_T_446_addr;
    GEN_13 <= T_406_2_T_446_en;
    if(T_406_2_T_437_en & T_406_2_T_437_mask) begin
      T_406_2[T_406_2_T_437_addr] <= T_406_2_T_437_data;
    end
    GEN_16 <= T_406_3_T_446_addr;
    GEN_18 <= T_406_3_T_446_en;
    if(T_406_3_T_437_en & T_406_3_T_437_mask) begin
      T_406_3[T_406_3_T_437_addr] <= T_406_3_T_437_data;
    end
    GEN_21 <= T_406_4_T_446_addr;
    GEN_23 <= T_406_4_T_446_en;
    if(T_406_4_T_437_en & T_406_4_T_437_mask) begin
      T_406_4[T_406_4_T_437_addr] <= T_406_4_T_437_data;
    end
    GEN_26 <= T_406_5_T_446_addr;
    GEN_29 <= T_406_5_T_446_en;
    if(T_406_5_T_437_en & T_406_5_T_437_mask) begin
      T_406_5[T_406_5_T_437_addr] <= T_406_5_T_437_data;
    end
    GEN_35 <= T_406_6_T_446_addr;
    GEN_39 <= T_406_6_T_446_en;
    if(T_406_6_T_437_en & T_406_6_T_437_mask) begin
      T_406_6[T_406_6_T_437_addr] <= T_406_6_T_437_data;
    end
    GEN_44 <= T_406_7_T_446_addr;
    GEN_46 <= T_406_7_T_446_en;
    if(T_406_7_T_437_en & T_406_7_T_437_mask) begin
      T_406_7[T_406_7_T_437_addr] <= T_406_7_T_437_data;
    end
  end
endmodule
module Arbiter_2(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [12:0] io_in_0_bits_addr,
  input   io_in_0_bits_write,
  input  [63:0] io_in_0_bits_wdata,
  input  [7:0] io_in_0_bits_wmask,
  input   io_in_0_bits_way_en,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [12:0] io_in_1_bits_addr,
  input   io_in_1_bits_write,
  input  [63:0] io_in_1_bits_wdata,
  input  [7:0] io_in_1_bits_wmask,
  input   io_in_1_bits_way_en,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [12:0] io_in_2_bits_addr,
  input   io_in_2_bits_write,
  input  [63:0] io_in_2_bits_wdata,
  input  [7:0] io_in_2_bits_wmask,
  input   io_in_2_bits_way_en,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [12:0] io_in_3_bits_addr,
  input   io_in_3_bits_write,
  input  [63:0] io_in_3_bits_wdata,
  input  [7:0] io_in_3_bits_wmask,
  input   io_in_3_bits_way_en,
  input   io_out_ready,
  output  io_out_valid,
  output [12:0] io_out_bits_addr,
  output  io_out_bits_write,
  output [63:0] io_out_bits_wdata,
  output [7:0] io_out_bits_wmask,
  output  io_out_bits_way_en,
  output [1:0] io_chosen
);
  wire [1:0] GEN_0;
  wire [12:0] GEN_1;
  wire  GEN_2;
  wire [63:0] GEN_3;
  wire [7:0] GEN_4;
  wire  GEN_5;
  wire [1:0] GEN_6;
  wire [12:0] GEN_7;
  wire  GEN_8;
  wire [63:0] GEN_9;
  wire [7:0] GEN_10;
  wire  GEN_11;
  wire [1:0] GEN_12;
  wire [12:0] GEN_13;
  wire  GEN_14;
  wire [63:0] GEN_15;
  wire [7:0] GEN_16;
  wire  GEN_17;
  wire  T_2025;
  wire  T_2026;
  wire  T_2028;
  wire  T_2030;
  wire  T_2032;
  wire  T_2034;
  wire  T_2035;
  wire  T_2036;
  wire  T_2038;
  wire  T_2039;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_2034;
  assign io_in_2_ready = T_2035;
  assign io_in_3_ready = T_2036;
  assign io_out_valid = T_2039;
  assign io_out_bits_addr = GEN_13;
  assign io_out_bits_write = GEN_14;
  assign io_out_bits_wdata = GEN_15;
  assign io_out_bits_wmask = GEN_16;
  assign io_out_bits_way_en = GEN_17;
  assign io_chosen = GEN_12;
  assign GEN_0 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_1 = io_in_2_valid ? io_in_2_bits_addr : io_in_3_bits_addr;
  assign GEN_2 = io_in_2_valid ? io_in_2_bits_write : io_in_3_bits_write;
  assign GEN_3 = io_in_2_valid ? io_in_2_bits_wdata : io_in_3_bits_wdata;
  assign GEN_4 = io_in_2_valid ? io_in_2_bits_wmask : io_in_3_bits_wmask;
  assign GEN_5 = io_in_2_valid ? io_in_2_bits_way_en : io_in_3_bits_way_en;
  assign GEN_6 = io_in_1_valid ? 2'h1 : GEN_0;
  assign GEN_7 = io_in_1_valid ? io_in_1_bits_addr : GEN_1;
  assign GEN_8 = io_in_1_valid ? io_in_1_bits_write : GEN_2;
  assign GEN_9 = io_in_1_valid ? io_in_1_bits_wdata : GEN_3;
  assign GEN_10 = io_in_1_valid ? io_in_1_bits_wmask : GEN_4;
  assign GEN_11 = io_in_1_valid ? io_in_1_bits_way_en : GEN_5;
  assign GEN_12 = io_in_0_valid ? 2'h0 : GEN_6;
  assign GEN_13 = io_in_0_valid ? io_in_0_bits_addr : GEN_7;
  assign GEN_14 = io_in_0_valid ? io_in_0_bits_write : GEN_8;
  assign GEN_15 = io_in_0_valid ? io_in_0_bits_wdata : GEN_9;
  assign GEN_16 = io_in_0_valid ? io_in_0_bits_wmask : GEN_10;
  assign GEN_17 = io_in_0_valid ? io_in_0_bits_way_en : GEN_11;
  assign T_2025 = io_in_0_valid | io_in_1_valid;
  assign T_2026 = T_2025 | io_in_2_valid;
  assign T_2028 = io_in_0_valid == 1'h0;
  assign T_2030 = T_2025 == 1'h0;
  assign T_2032 = T_2026 == 1'h0;
  assign T_2034 = T_2028 & io_out_ready;
  assign T_2035 = T_2030 & io_out_ready;
  assign T_2036 = T_2032 & io_out_ready;
  assign T_2038 = T_2032 == 1'h0;
  assign T_2039 = T_2038 | io_in_3_valid;
endmodule
module DCache(
  input   clk,
  input   reset,
  output  io_cpu_req_ready,
  input   io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_addr,
  input  [8:0] io_cpu_req_bits_tag,
  input  [4:0] io_cpu_req_bits_cmd,
  input  [2:0] io_cpu_req_bits_typ,
  input   io_cpu_req_bits_phys,
  input  [31:0] io_cpu_req_bits_data,
  input   io_cpu_s1_kill,
  input  [31:0] io_cpu_s1_data,
  output  io_cpu_s2_nack,
  output  io_cpu_resp_valid,
  output [31:0] io_cpu_resp_bits_addr,
  output [8:0] io_cpu_resp_bits_tag,
  output [4:0] io_cpu_resp_bits_cmd,
  output [2:0] io_cpu_resp_bits_typ,
  output [31:0] io_cpu_resp_bits_data,
  output  io_cpu_resp_bits_replay,
  output  io_cpu_resp_bits_has_data,
  output [31:0] io_cpu_resp_bits_data_word_bypass,
  output [31:0] io_cpu_resp_bits_store_data,
  output  io_cpu_replay_next,
  output  io_cpu_xcpt_ma_ld,
  output  io_cpu_xcpt_ma_st,
  output  io_cpu_xcpt_pf_ld,
  output  io_cpu_xcpt_pf_st,
  input   io_cpu_invalidate_lr,
  output  io_cpu_ordered,
  input   io_ptw_req_ready,
  output  io_ptw_req_valid,
  output [1:0] io_ptw_req_bits_prv,
  output  io_ptw_req_bits_pum,
  output  io_ptw_req_bits_mxr,
  output [19:0] io_ptw_req_bits_addr,
  output  io_ptw_req_bits_store,
  output  io_ptw_req_bits_fetch,
  input   io_ptw_resp_valid,
  input  [15:0] io_ptw_resp_bits_pte_reserved_for_hardware,
  input  [37:0] io_ptw_resp_bits_pte_ppn,
  input  [1:0] io_ptw_resp_bits_pte_reserved_for_software,
  input   io_ptw_resp_bits_pte_d,
  input   io_ptw_resp_bits_pte_a,
  input   io_ptw_resp_bits_pte_g,
  input   io_ptw_resp_bits_pte_u,
  input   io_ptw_resp_bits_pte_x,
  input   io_ptw_resp_bits_pte_w,
  input   io_ptw_resp_bits_pte_r,
  input   io_ptw_resp_bits_pte_v,
  input  [6:0] io_ptw_ptbr_asid,
  input  [21:0] io_ptw_ptbr_ppn,
  input   io_ptw_invalidate,
  input   io_ptw_status_debug,
  input  [1:0] io_ptw_status_prv,
  input   io_ptw_status_sd,
  input  [30:0] io_ptw_status_zero3,
  input   io_ptw_status_sd_rv32,
  input  [1:0] io_ptw_status_zero2,
  input  [4:0] io_ptw_status_vm,
  input  [3:0] io_ptw_status_zero1,
  input   io_ptw_status_mxr,
  input   io_ptw_status_pum,
  input   io_ptw_status_mprv,
  input  [1:0] io_ptw_status_xs,
  input  [1:0] io_ptw_status_fs,
  input  [1:0] io_ptw_status_mpp,
  input  [1:0] io_ptw_status_hpp,
  input   io_ptw_status_spp,
  input   io_ptw_status_mpie,
  input   io_ptw_status_hpie,
  input   io_ptw_status_spie,
  input   io_ptw_status_upie,
  input   io_ptw_status_mie,
  input   io_ptw_status_hie,
  input   io_ptw_status_sie,
  input   io_ptw_status_uie,
  input   io_mem_acquire_ready,
  output  io_mem_acquire_valid,
  output [25:0] io_mem_acquire_bits_addr_block,
  output  io_mem_acquire_bits_client_xact_id,
  output [2:0] io_mem_acquire_bits_addr_beat,
  output  io_mem_acquire_bits_is_builtin_type,
  output [2:0] io_mem_acquire_bits_a_type,
  output [11:0] io_mem_acquire_bits_union,
  output [63:0] io_mem_acquire_bits_data,
  output  io_mem_probe_ready,
  input   io_mem_probe_valid,
  input  [25:0] io_mem_probe_bits_addr_block,
  input  [1:0] io_mem_probe_bits_p_type,
  input   io_mem_release_ready,
  output  io_mem_release_valid,
  output [2:0] io_mem_release_bits_addr_beat,
  output [25:0] io_mem_release_bits_addr_block,
  output  io_mem_release_bits_client_xact_id,
  output  io_mem_release_bits_voluntary,
  output [2:0] io_mem_release_bits_r_type,
  output [63:0] io_mem_release_bits_data,
  output  io_mem_grant_ready,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input   io_mem_grant_bits_client_xact_id,
  input  [1:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data,
  input   io_mem_grant_bits_manager_id,
  input   io_mem_finish_ready,
  output  io_mem_finish_valid,
  output [1:0] io_mem_finish_bits_manager_xact_id,
  output  io_mem_finish_bits_manager_id
);
  wire  fq_clk;
  wire  fq_reset;
  wire  fq_io_enq_ready;
  wire  fq_io_enq_valid;
  wire [1:0] fq_io_enq_bits_manager_xact_id;
  wire  fq_io_enq_bits_manager_id;
  wire  fq_io_deq_ready;
  wire  fq_io_deq_valid;
  wire [1:0] fq_io_deq_bits_manager_xact_id;
  wire  fq_io_deq_bits_manager_id;
  wire  fq_io_count;
  wire  T_1924;
  reg [15:0] T_1927;
  reg [31:0] GEN_48;
  wire  T_1928;
  wire  T_1929;
  wire  T_1930;
  wire  T_1931;
  wire  T_1932;
  wire  T_1933;
  wire  T_1934;
  wire [14:0] T_1935;
  wire [15:0] T_1936;
  wire [15:0] GEN_2;
  wire  meta_clk;
  wire  meta_reset;
  wire  meta_io_read_ready;
  wire  meta_io_read_valid;
  wire [6:0] meta_io_read_bits_idx;
  wire  meta_io_read_bits_way_en;
  wire  meta_io_write_ready;
  wire  meta_io_write_valid;
  wire [6:0] meta_io_write_bits_idx;
  wire  meta_io_write_bits_way_en;
  wire [18:0] meta_io_write_bits_data_tag;
  wire [1:0] meta_io_write_bits_data_coh_state;
  wire [18:0] meta_io_resp_0_tag;
  wire [1:0] meta_io_resp_0_coh_state;
  wire  metaReadArb_clk;
  wire  metaReadArb_reset;
  wire  metaReadArb_io_in_0_ready;
  wire  metaReadArb_io_in_0_valid;
  wire [6:0] metaReadArb_io_in_0_bits_idx;
  wire  metaReadArb_io_in_0_bits_way_en;
  wire  metaReadArb_io_in_1_ready;
  wire  metaReadArb_io_in_1_valid;
  wire [6:0] metaReadArb_io_in_1_bits_idx;
  wire  metaReadArb_io_in_1_bits_way_en;
  wire  metaReadArb_io_in_2_ready;
  wire  metaReadArb_io_in_2_valid;
  wire [6:0] metaReadArb_io_in_2_bits_idx;
  wire  metaReadArb_io_in_2_bits_way_en;
  wire  metaReadArb_io_out_ready;
  wire  metaReadArb_io_out_valid;
  wire [6:0] metaReadArb_io_out_bits_idx;
  wire  metaReadArb_io_out_bits_way_en;
  wire [1:0] metaReadArb_io_chosen;
  wire  metaWriteArb_clk;
  wire  metaWriteArb_reset;
  wire  metaWriteArb_io_in_0_ready;
  wire  metaWriteArb_io_in_0_valid;
  wire [6:0] metaWriteArb_io_in_0_bits_idx;
  wire  metaWriteArb_io_in_0_bits_way_en;
  wire [18:0] metaWriteArb_io_in_0_bits_data_tag;
  wire [1:0] metaWriteArb_io_in_0_bits_data_coh_state;
  wire  metaWriteArb_io_in_1_ready;
  wire  metaWriteArb_io_in_1_valid;
  wire [6:0] metaWriteArb_io_in_1_bits_idx;
  wire  metaWriteArb_io_in_1_bits_way_en;
  wire [18:0] metaWriteArb_io_in_1_bits_data_tag;
  wire [1:0] metaWriteArb_io_in_1_bits_data_coh_state;
  wire  metaWriteArb_io_in_2_ready;
  wire  metaWriteArb_io_in_2_valid;
  wire [6:0] metaWriteArb_io_in_2_bits_idx;
  wire  metaWriteArb_io_in_2_bits_way_en;
  wire [18:0] metaWriteArb_io_in_2_bits_data_tag;
  wire [1:0] metaWriteArb_io_in_2_bits_data_coh_state;
  wire  metaWriteArb_io_out_ready;
  wire  metaWriteArb_io_out_valid;
  wire [6:0] metaWriteArb_io_out_bits_idx;
  wire  metaWriteArb_io_out_bits_way_en;
  wire [18:0] metaWriteArb_io_out_bits_data_tag;
  wire [1:0] metaWriteArb_io_out_bits_data_coh_state;
  wire [1:0] metaWriteArb_io_chosen;
  wire  data_clk;
  wire  data_reset;
  wire  data_io_req_valid;
  wire [12:0] data_io_req_bits_addr;
  wire  data_io_req_bits_write;
  wire [63:0] data_io_req_bits_wdata;
  wire [7:0] data_io_req_bits_wmask;
  wire  data_io_req_bits_way_en;
  wire [63:0] data_io_resp_0;
  wire  dataArb_clk;
  wire  dataArb_reset;
  wire  dataArb_io_in_0_ready;
  wire  dataArb_io_in_0_valid;
  wire [12:0] dataArb_io_in_0_bits_addr;
  wire  dataArb_io_in_0_bits_write;
  wire [63:0] dataArb_io_in_0_bits_wdata;
  wire [7:0] dataArb_io_in_0_bits_wmask;
  wire  dataArb_io_in_0_bits_way_en;
  wire  dataArb_io_in_1_ready;
  wire  dataArb_io_in_1_valid;
  wire [12:0] dataArb_io_in_1_bits_addr;
  wire  dataArb_io_in_1_bits_write;
  wire [63:0] dataArb_io_in_1_bits_wdata;
  wire [7:0] dataArb_io_in_1_bits_wmask;
  wire  dataArb_io_in_1_bits_way_en;
  wire  dataArb_io_in_2_ready;
  wire  dataArb_io_in_2_valid;
  wire [12:0] dataArb_io_in_2_bits_addr;
  wire  dataArb_io_in_2_bits_write;
  wire [63:0] dataArb_io_in_2_bits_wdata;
  wire [7:0] dataArb_io_in_2_bits_wmask;
  wire  dataArb_io_in_2_bits_way_en;
  wire  dataArb_io_in_3_ready;
  wire  dataArb_io_in_3_valid;
  wire [12:0] dataArb_io_in_3_bits_addr;
  wire  dataArb_io_in_3_bits_write;
  wire [63:0] dataArb_io_in_3_bits_wdata;
  wire [7:0] dataArb_io_in_3_bits_wmask;
  wire  dataArb_io_in_3_bits_way_en;
  wire  dataArb_io_out_ready;
  wire  dataArb_io_out_valid;
  wire [12:0] dataArb_io_out_bits_addr;
  wire  dataArb_io_out_bits_write;
  wire [63:0] dataArb_io_out_bits_wdata;
  wire [7:0] dataArb_io_out_bits_wmask;
  wire  dataArb_io_out_bits_way_en;
  wire [1:0] dataArb_io_chosen;
  wire  T_2218;
  reg  s1_valid;
  reg [31:0] GEN_49;
  wire  T_2220;
  reg  s1_probe;
  reg [31:0] GEN_50;
  reg [25:0] probe_bits_addr_block;
  reg [31:0] GEN_51;
  reg [1:0] probe_bits_p_type;
  reg [31:0] GEN_52;
  wire [25:0] GEN_3;
  wire [1:0] GEN_4;
  wire  s1_nack;
  wire  T_2247;
  wire  s1_valid_masked;
  wire  T_2249;
  wire  s1_valid_not_nacked;
  reg [31:0] s1_req_addr;
  reg [31:0] GEN_53;
  reg [8:0] s1_req_tag;
  reg [31:0] GEN_75;
  reg [4:0] s1_req_cmd;
  reg [31:0] GEN_88;
  reg [2:0] s1_req_typ;
  reg [31:0] GEN_89;
  reg  s1_req_phys;
  reg [31:0] GEN_93;
  reg [31:0] s1_req_data;
  reg [31:0] GEN_97;
  wire [18:0] T_2316;
  wire [5:0] T_2317;
  wire [25:0] T_2318;
  wire [31:0] T_2319;
  wire [31:0] GEN_5;
  wire [8:0] GEN_6;
  wire [4:0] GEN_7;
  wire [2:0] GEN_8;
  wire  GEN_9;
  wire [31:0] GEN_10;
  wire  T_2320;
  wire  T_2321;
  wire  T_2322;
  wire  T_2323;
  wire  T_2324;
  wire  T_2325;
  wire  T_2326;
  wire  T_2327;
  wire  s1_read;
  wire  T_2328;
  wire  T_2330;
  wire  s1_write;
  wire  s1_readwrite;
  reg  s1_flush_valid;
  reg [31:0] GEN_98;
  reg  grant_wait;
  reg [31:0] GEN_102;
  reg  release_ack_wait;
  reg [31:0] GEN_110;
  reg [2:0] release_state;
  reg [31:0] GEN_119;
  wire  pstore1_valid;
  reg  pstore2_valid;
  reg [31:0] GEN_133;
  wire  T_2340;
  wire  T_2341;
  wire  inWriteback;
  wire [1:0] releaseWay;
  wire  T_2343;
  wire  T_2345;
  wire  T_2346;
  wire  T_2349;
  wire  T_2350;
  wire  T_2351;
  wire  T_2352;
  wire  T_2353;
  wire  T_2354;
  wire  T_2355;
  wire  T_2356;
  wire  T_2357;
  wire  T_2358;
  wire  T_2359;
  wire  T_2364;
  wire  T_2374;
  wire  GEN_11;
  wire [6:0] T_2376;
  wire  T_2380;
  wire  GEN_12;
  wire  tlb_clk;
  wire  tlb_reset;
  wire  tlb_io_req_ready;
  wire  tlb_io_req_valid;
  wire [19:0] tlb_io_req_bits_vpn;
  wire  tlb_io_req_bits_passthrough;
  wire  tlb_io_req_bits_instruction;
  wire  tlb_io_req_bits_store;
  wire  tlb_io_resp_miss;
  wire [19:0] tlb_io_resp_ppn;
  wire  tlb_io_resp_xcpt_ld;
  wire  tlb_io_resp_xcpt_st;
  wire  tlb_io_resp_xcpt_if;
  wire  tlb_io_resp_cacheable;
  wire  tlb_io_ptw_req_ready;
  wire  tlb_io_ptw_req_valid;
  wire [1:0] tlb_io_ptw_req_bits_prv;
  wire  tlb_io_ptw_req_bits_pum;
  wire  tlb_io_ptw_req_bits_mxr;
  wire [19:0] tlb_io_ptw_req_bits_addr;
  wire  tlb_io_ptw_req_bits_store;
  wire  tlb_io_ptw_req_bits_fetch;
  wire  tlb_io_ptw_resp_valid;
  wire [15:0] tlb_io_ptw_resp_bits_pte_reserved_for_hardware;
  wire [37:0] tlb_io_ptw_resp_bits_pte_ppn;
  wire [1:0] tlb_io_ptw_resp_bits_pte_reserved_for_software;
  wire  tlb_io_ptw_resp_bits_pte_d;
  wire  tlb_io_ptw_resp_bits_pte_a;
  wire  tlb_io_ptw_resp_bits_pte_g;
  wire  tlb_io_ptw_resp_bits_pte_u;
  wire  tlb_io_ptw_resp_bits_pte_x;
  wire  tlb_io_ptw_resp_bits_pte_w;
  wire  tlb_io_ptw_resp_bits_pte_r;
  wire  tlb_io_ptw_resp_bits_pte_v;
  wire [6:0] tlb_io_ptw_ptbr_asid;
  wire [21:0] tlb_io_ptw_ptbr_ppn;
  wire  tlb_io_ptw_invalidate;
  wire  tlb_io_ptw_status_debug;
  wire [1:0] tlb_io_ptw_status_prv;
  wire  tlb_io_ptw_status_sd;
  wire [30:0] tlb_io_ptw_status_zero3;
  wire  tlb_io_ptw_status_sd_rv32;
  wire [1:0] tlb_io_ptw_status_zero2;
  wire [4:0] tlb_io_ptw_status_vm;
  wire [3:0] tlb_io_ptw_status_zero1;
  wire  tlb_io_ptw_status_mxr;
  wire  tlb_io_ptw_status_pum;
  wire  tlb_io_ptw_status_mprv;
  wire [1:0] tlb_io_ptw_status_xs;
  wire [1:0] tlb_io_ptw_status_fs;
  wire [1:0] tlb_io_ptw_status_mpp;
  wire [1:0] tlb_io_ptw_status_hpp;
  wire  tlb_io_ptw_status_spp;
  wire  tlb_io_ptw_status_mpie;
  wire  tlb_io_ptw_status_hpie;
  wire  tlb_io_ptw_status_spie;
  wire  tlb_io_ptw_status_upie;
  wire  tlb_io_ptw_status_mie;
  wire  tlb_io_ptw_status_hie;
  wire  tlb_io_ptw_status_sie;
  wire  tlb_io_ptw_status_uie;
  wire  T_2382;
  wire [19:0] T_2383;
  wire  T_2386;
  wire  T_2388;
  wire  T_2389;
  wire  GEN_13;
  wire  T_2391;
  wire  T_2392;
  wire [11:0] T_2394;
  wire [31:0] s1_paddr;
  wire [18:0] T_2395;
  wire [18:0] T_2396;
  wire [18:0] s1_tag;
  wire  T_2397;
  wire  T_2398;
  wire  s1_hit_way;
  wire [1:0] T_2422_state;
  wire [1:0] T_2446;
  wire [1:0] s1_hit_state_state;
  wire  s1_victim_way;
  reg  s2_valid;
  reg [31:0] GEN_134;
  reg  s2_probe;
  reg [31:0] GEN_135;
  wire  T_2496;
  wire  T_2497;
  wire  releaseInFlight;
  reg  T_2500;
  reg [31:0] GEN_136;
  wire  s2_valid_masked;
  reg [31:0] s2_req_addr;
  reg [31:0] GEN_137;
  reg [8:0] s2_req_tag;
  reg [31:0] GEN_138;
  reg [4:0] s2_req_cmd;
  reg [31:0] GEN_139;
  reg [2:0] s2_req_typ;
  reg [31:0] GEN_140;
  reg  s2_req_phys;
  reg [31:0] GEN_141;
  reg [31:0] s2_req_data;
  reg [31:0] GEN_142;
  reg  s2_uncached;
  reg [31:0] GEN_143;
  wire  T_2568;
  wire  T_2570;
  wire [31:0] GEN_15;
  wire [8:0] GEN_16;
  wire [4:0] GEN_17;
  wire [2:0] GEN_18;
  wire  GEN_19;
  wire [31:0] GEN_20;
  wire  GEN_21;
  wire  T_2571;
  wire  T_2572;
  wire  T_2573;
  wire  T_2574;
  wire  T_2575;
  wire  T_2576;
  wire  T_2577;
  wire  T_2578;
  wire  s2_read;
  wire  T_2579;
  wire  T_2581;
  wire  s2_write;
  wire  s2_readwrite;
  reg  s2_flush_valid;
  reg [31:0] GEN_144;
  wire  T_2585;
  reg [63:0] s2_data;
  reg [63:0] GEN_145;
  wire [63:0] GEN_22;
  reg  s2_probe_way;
  reg [31:0] GEN_146;
  wire  GEN_23;
  reg [1:0] s2_probe_state_state;
  reg [31:0] GEN_147;
  wire [1:0] GEN_24;
  reg  s2_hit_way;
  reg [31:0] GEN_148;
  wire  GEN_25;
  reg [1:0] s2_hit_state_state;
  reg [31:0] GEN_149;
  wire [1:0] GEN_26;
  wire  T_2635;
  wire  T_2636;
  wire  T_2638;
  wire  T_2639;
  wire  T_2640;
  wire  T_2641;
  wire  s2_hit;
  wire  T_2645;
  wire  s2_valid_hit;
  wire  T_2648;
  wire  T_2649;
  wire  T_2650;
  wire  T_2652;
  wire  T_2653;
  wire  T_2655;
  wire  s2_valid_miss;
  wire  T_2657;
  wire  s2_valid_cached_miss;
  wire  s2_victimize;
  wire  s2_valid_uncached;
  wire  T_2658;
  wire  T_2660;
  wire  T_2661;
  reg  T_2663;
  reg [31:0] GEN_150;
  wire  GEN_27;
  wire [1:0] T_2665;
  wire [1:0] s2_victim_way;
  reg [18:0] s2_victim_tag;
  reg [31:0] GEN_151;
  wire [18:0] GEN_0;
  wire [18:0] GEN_28;
  wire [18:0] GEN_29;
  reg [1:0] T_2839_state;
  reg [31:0] GEN_152;
  wire [1:0] GEN_1;
  wire [1:0] GEN_30;
  wire [1:0] GEN_31;
  wire [1:0] s2_victim_state_state;
  wire  s2_victim_dirty;
  wire  T_2883;
  wire  T_2884;
  wire  T_2885;
  wire  T_2887;
  wire  T_2888;
  wire  GEN_32;
  wire [1:0] T_2894;
  wire [3:0] T_2896;
  wire [4:0] T_2898;
  wire [3:0] T_2899;
  wire [1:0] T_2900;
  wire [31:0] GEN_123;
  wire [31:0] T_2901;
  wire  misaligned;
  wire  T_2903;
  wire  T_2904;
  wire  T_2905;
  wire  T_2906;
  wire  T_2907;
  wire  T_2908;
  wire  T_2909;
  reg  T_2910;
  reg [31:0] GEN_153;
  wire  T_2911;
  wire  T_2913;
  wire  T_2914;
  wire  T_2916;
  reg [4:0] lrscCount;
  reg [31:0] GEN_154;
  wire  lrscValid;
  reg [25:0] lrscAddr;
  reg [31:0] GEN_155;
  wire [5:0] T_2933;
  wire [4:0] T_2934;
  wire [4:0] GEN_35;
  wire [4:0] GEN_36;
  wire  T_2938;
  reg [4:0] pstore1_cmd;
  reg [31:0] GEN_156;
  wire [4:0] GEN_37;
  reg [2:0] pstore1_typ;
  reg [31:0] GEN_157;
  wire [2:0] GEN_38;
  reg [31:0] pstore1_addr;
  reg [31:0] GEN_158;
  wire [31:0] GEN_39;
  reg [31:0] pstore1_data;
  reg [31:0] GEN_159;
  wire [31:0] GEN_40;
  reg  pstore1_way;
  reg [31:0] GEN_160;
  wire  GEN_41;
  wire [1:0] T_2943;
  wire  T_2945;
  wire [7:0] T_2946;
  wire [15:0] T_2947;
  wire [31:0] T_2948;
  wire  T_2950;
  wire [15:0] T_2951;
  wire [31:0] T_2952;
  wire [31:0] T_2953;
  wire [31:0] T_2954;
  wire [31:0] pstore1_storegen_data;
  wire  pstore_drain_opportunistic;
  wire  pstore_drain_on_miss;
  wire  T_2985;
  wire  T_2986;
  wire  T_2987;
  reg  T_2992;
  reg [31:0] GEN_161;
  wire  T_2994;
  wire  T_2996;
  wire  T_2997;
  wire  T_2998;
  wire  T_3000;
  wire  T_3001;
  wire  T_3002;
  wire  T_3004;
  wire  T_3005;
  wire  T_3007;
  wire  advance_pstore1;
  wire  T_3010;
  wire  T_3011;
  reg [31:0] pstore2_addr;
  reg [31:0] GEN_162;
  wire [31:0] GEN_42;
  reg  pstore2_way;
  reg [31:0] GEN_163;
  wire  GEN_43;
  reg [31:0] pstore2_storegen_data;
  reg [31:0] GEN_164;
  wire [31:0] GEN_44;
  wire  T_3013;
  wire  T_3017;
  wire  T_3021;
  wire  T_3024;
  wire [1:0] T_3025;
  wire  T_3026;
  wire [1:0] T_3028;
  wire  T_3030;
  wire [1:0] T_3033;
  wire [1:0] T_3034;
  wire [1:0] T_3037;
  wire [3:0] T_3038;
  reg [3:0] pstore2_storegen_mask;
  reg [31:0] GEN_165;
  wire [3:0] GEN_45;
  wire [31:0] T_3040;
  wire  T_3041;
  wire [31:0] T_3042;
  wire [63:0] T_3043;
  wire  T_3045;
  wire [2:0] GEN_124;
  wire [2:0] pstore_mask_shift;
  wire [3:0] T_3073;
  wire [10:0] GEN_125;
  wire [10:0] T_3074;
  wire [10:0] s1_idx;
  wire [10:0] T_3075;
  wire  T_3076;
  wire  T_3077;
  wire [10:0] T_3078;
  wire  T_3079;
  wire  T_3080;
  wire  T_3081;
  wire  s1_raw_hazard;
  wire  T_3082;
  wire  GEN_46;
  wire [1:0] T_3091;
  wire [1:0] s2_new_hit_state_state;
  wire  T_3135;
  wire  T_3137;
  wire  T_3138;
  wire  T_3140;
  wire  T_3141;
  wire  T_3142;
  wire [6:0] T_3143;
  wire [1:0] T_3167_state;
  wire [1:0] T_3189_state;
  wire [18:0] T_3211;
  wire [25:0] T_3213;
  wire [5:0] T_3228;
  wire [25:0] cachedGetMessage_addr_block;
  wire  cachedGetMessage_client_xact_id;
  wire [2:0] cachedGetMessage_addr_beat;
  wire  cachedGetMessage_is_builtin_type;
  wire [2:0] cachedGetMessage_a_type;
  wire [11:0] cachedGetMessage_union;
  wire [63:0] cachedGetMessage_data;
  wire [2:0] T_3288;
  wire [2:0] T_3289;
  wire [5:0] T_3330;
  wire [11:0] T_3331;
  wire [25:0] uncachedGetMessage_addr_block;
  wire  uncachedGetMessage_client_xact_id;
  wire [2:0] uncachedGetMessage_addr_beat;
  wire  uncachedGetMessage_is_builtin_type;
  wire [2:0] uncachedGetMessage_a_type;
  wire [11:0] uncachedGetMessage_union;
  wire [63:0] uncachedGetMessage_data;
  wire  uncachedPutOffset;
  wire [63:0] T_3430;
  wire [2:0] GEN_126;
  wire [2:0] T_3458;
  wire [10:0] GEN_127;
  wire [10:0] T_3459;
  wire [7:0] T_3496;
  wire [8:0] T_3506;
  wire [11:0] T_3526;
  wire [25:0] uncachedPutMessage_addr_block;
  wire  uncachedPutMessage_client_xact_id;
  wire [2:0] uncachedPutMessage_addr_beat;
  wire  uncachedPutMessage_is_builtin_type;
  wire [2:0] uncachedPutMessage_a_type;
  wire [11:0] uncachedPutMessage_union;
  wire [63:0] uncachedPutMessage_data;
  wire [11:0] T_3642;
  wire [25:0] uncachedPutAtomicMessage_addr_block;
  wire  uncachedPutAtomicMessage_client_xact_id;
  wire [2:0] uncachedPutAtomicMessage_addr_beat;
  wire  uncachedPutAtomicMessage_is_builtin_type;
  wire [2:0] uncachedPutAtomicMessage_a_type;
  wire [11:0] uncachedPutAtomicMessage_union;
  wire [63:0] uncachedPutAtomicMessage_data;
  wire  T_3729;
  wire  T_3730;
  wire  T_3731;
  wire  T_3733;
  wire  T_3736;
  wire  T_3737;
  wire  T_3738;
  wire  T_3740;
  wire [25:0] GEN_54;
  wire  GEN_55;
  wire [2:0] GEN_56;
  wire  GEN_57;
  wire [2:0] GEN_58;
  wire [11:0] GEN_59;
  wire [63:0] GEN_60;
  wire [25:0] GEN_61;
  wire  GEN_62;
  wire [2:0] GEN_63;
  wire  GEN_64;
  wire [2:0] GEN_65;
  wire [11:0] GEN_66;
  wire [63:0] GEN_67;
  wire  T_3741;
  wire  GEN_68;
  wire [2:0] T_3750_0;
  wire [3:0] GEN_128;
  wire  T_3752;
  wire  T_3753;
  wire  T_3754;
  wire  grantIsVoluntary;
  wire  T_3758;
  wire  T_3760;
  wire  grantIsUncached;
  wire  T_3761;
  wire  T_3762;
  wire  T_3763;
  wire  T_3765;
  wire [63:0] GEN_69;
  wire  GEN_70;
  wire [63:0] GEN_71;
  wire  GEN_72;
  wire  T_3767;
  wire  T_3768;
  reg [2:0] refillCount;
  reg [31:0] GEN_166;
  wire  T_3771;
  wire [3:0] T_3773;
  wire [2:0] T_3774;
  wire [2:0] GEN_73;
  wire  refillDone;
  wire  grantDone;
  wire  T_3776;
  wire  GEN_74;
  wire  T_3778;
  wire  T_3781;
  wire  T_3782;
  wire  T_3783;
  wire  T_3785;
  wire [28:0] T_3788;
  wire [31:0] GEN_129;
  wire [31:0] T_3789;
  wire  T_3793;
  wire  T_3794;
  wire  T_3795;
  wire  T_3797;
  wire [1:0] T_3806;
  wire [1:0] T_3807;
  wire [1:0] T_3830_state;
  wire  T_3863;
  wire  T_3866;
  wire  T_3867;
  wire [1:0] T_3891_manager_xact_id;
  wire  T_3891_manager_id;
  wire  T_3914;
  wire  T_3916;
  wire  T_3918;
  wire  T_3921;
  wire  T_3922;
  wire  T_3925;
  wire  T_3927;
  wire  T_3928;
  wire  T_3930;
  wire  T_3931;
  wire  T_3932;
  wire  T_3935;
  wire  T_3936;
  reg [2:0] writebackCount;
  reg [31:0] GEN_167;
  wire  T_3939;
  wire [3:0] T_3941;
  wire [2:0] T_3942;
  wire [2:0] GEN_76;
  wire  writebackDone;
  wire  T_3945;
  wire  T_3946;
  wire  releaseDone;
  wire  T_3948;
  wire  releaseRejected;
  wire  T_3949;
  reg  s1_release_data_valid;
  reg [31:0] GEN_168;
  wire  T_3951;
  wire  T_3952;
  reg  s2_release_data_valid;
  reg [31:0] GEN_169;
  wire [3:0] T_3954;
  wire [1:0] T_3957;
  wire [1:0] GEN_130;
  wire [2:0] T_3958;
  wire [1:0] T_3959;
  wire [1:0] T_3960;
  wire [3:0] GEN_131;
  wire [4:0] T_3961;
  wire [3:0] releaseDataBeat;
  wire [1:0] T_3985_state;
  wire  T_4010;
  wire [2:0] T_4011;
  wire  T_4040;
  wire [2:0] T_4041;
  wire  T_4042;
  wire [2:0] T_4043;
  wire  T_4044;
  wire [2:0] T_4045;
  wire [2:0] T_4074_addr_beat;
  wire [25:0] T_4074_addr_block;
  wire  T_4074_client_xact_id;
  wire  T_4074_voluntary;
  wire [2:0] T_4074_r_type;
  wire [63:0] T_4074_data;
  wire [2:0] T_4107;
  wire [2:0] voluntaryReleaseMessage_addr_beat;
  wire [25:0] voluntaryReleaseMessage_addr_block;
  wire  voluntaryReleaseMessage_client_xact_id;
  wire  voluntaryReleaseMessage_voluntary;
  wire [2:0] voluntaryReleaseMessage_r_type;
  wire [63:0] voluntaryReleaseMessage_data;
  wire [1:0] voluntaryNewCoh_state;
  wire  T_4221;
  wire [2:0] T_4222;
  wire [2:0] T_4252;
  wire [2:0] T_4254;
  wire [2:0] T_4256;
  wire [2:0] probeResponseMessage_addr_beat;
  wire [25:0] probeResponseMessage_addr_block;
  wire  probeResponseMessage_client_xact_id;
  wire  probeResponseMessage_voluntary;
  wire [2:0] probeResponseMessage_r_type;
  wire [63:0] probeResponseMessage_data;
  wire [1:0] T_4312;
  wire [1:0] T_4314;
  wire [1:0] T_4316;
  wire [1:0] probeNewCoh_state;
  wire [1:0] newCoh_state;
  wire  T_4381;
  wire  T_4385;
  wire  T_4387;
  wire [25:0] T_4389;
  wire [2:0] GEN_77;
  wire [25:0] GEN_78;
  wire [2:0] GEN_79;
  wire  T_4391;
  wire  T_4393;
  wire  T_4394;
  wire [2:0] GEN_80;
  wire  T_4398;
  wire  T_4399;
  wire  GEN_81;
  wire [2:0] GEN_82;
  wire [2:0] GEN_83;
  wire  GEN_84;
  wire [2:0] GEN_85;
  wire  T_4401;
  wire  T_4402;
  wire  T_4403;
  wire  GEN_86;
  wire  T_4407;
  wire [2:0] GEN_87;
  wire  GEN_90;
  wire  GEN_91;
  wire [2:0] GEN_92;
  wire [2:0] GEN_94;
  wire  T_4409;
  wire  T_4410;
  wire [2:0] GEN_95;
  wire  GEN_96;
  wire  GEN_99;
  wire  GEN_100;
  wire [2:0] GEN_101;
  wire [1:0] GEN_103;
  wire [1:0] GEN_104;
  wire [2:0] GEN_105;
  wire  GEN_106;
  wire  T_4414;
  wire  T_4415;
  wire  GEN_107;
  wire  T_4418;
  wire  T_4419;
  wire [2:0] T_4421;
  wire [28:0] T_4422;
  wire [31:0] GEN_132;
  wire [31:0] T_4423;
  wire  T_4427;
  wire  T_4428;
  wire [28:0] T_4430;
  wire [31:0] T_4431;
  wire [6:0] T_4432;
  wire [18:0] T_4436;
  wire  T_4437;
  wire [2:0] GEN_108;
  wire  T_4439;
  wire  T_4440;
  wire  T_4442;
  wire  T_4443;
  reg  doUncachedResp;
  reg [31:0] GEN_170;
  wire  T_4446;
  wire  T_4448;
  wire  GEN_109;
  wire [5:0] T_4452;
  wire [63:0] s2_data_word;
  wire [1:0] T_4453;
  wire [2:0] T_4454;
  wire  T_4456;
  wire  T_4457;
  wire [15:0] T_4458;
  wire [15:0] T_4459;
  wire [15:0] T_4460;
  wire  T_4466;
  wire  T_4468;
  wire  T_4469;
  wire [15:0] T_4473;
  wire [15:0] T_4475;
  wire [31:0] T_4476;
  wire  T_4477;
  wire [7:0] T_4478;
  wire [7:0] T_4479;
  wire [7:0] T_4480;
  wire  T_4486;
  wire  T_4488;
  wire  T_4489;
  wire [23:0] T_4493;
  wire [23:0] T_4494;
  wire [23:0] T_4495;
  wire [31:0] T_4496;
  wire  T_4498;
  wire  T_4499;
  wire  T_4501;
  wire  T_4502;
  wire  T_4504;
  reg  flushed;
  reg [31:0] GEN_171;
  reg  flushing;
  reg [31:0] GEN_172;
  reg [6:0] T_4508;
  reg [31:0] GEN_173;
  wire  GEN_111;
  wire  T_4511;
  wire  T_4512;
  wire  T_4514;
  wire  GEN_112;
  wire  GEN_113;
  wire  GEN_114;
  wire  T_4519;
  wire  T_4521;
  wire  T_4522;
  wire  T_4525;
  wire  T_4527;
  wire  T_4530;
  wire  T_4535;
  wire [7:0] T_4537;
  wire [6:0] T_4538;
  wire  GEN_115;
  wire [6:0] GEN_116;
  wire  GEN_117;
  wire  T_4541;
  wire  T_4544;
  wire  GEN_118;
  wire [6:0] GEN_120;
  wire  GEN_121;
  wire  GEN_122;
  reg [63:0] GEN_14;
  reg [63:0] GEN_174;
  reg [7:0] GEN_33;
  reg [31:0] GEN_175;
  reg [63:0] GEN_34;
  reg [63:0] GEN_176;
  reg [7:0] GEN_47;
  reg [31:0] GEN_177;
  FinishQueue fq (
    .clk(fq_clk),
    .reset(fq_reset),
    .io_enq_ready(fq_io_enq_ready),
    .io_enq_valid(fq_io_enq_valid),
    .io_enq_bits_manager_xact_id(fq_io_enq_bits_manager_xact_id),
    .io_enq_bits_manager_id(fq_io_enq_bits_manager_id),
    .io_deq_ready(fq_io_deq_ready),
    .io_deq_valid(fq_io_deq_valid),
    .io_deq_bits_manager_xact_id(fq_io_deq_bits_manager_xact_id),
    .io_deq_bits_manager_id(fq_io_deq_bits_manager_id),
    .io_count(fq_io_count)
  );
  MetadataArray meta (
    .clk(meta_clk),
    .reset(meta_reset),
    .io_read_ready(meta_io_read_ready),
    .io_read_valid(meta_io_read_valid),
    .io_read_bits_idx(meta_io_read_bits_idx),
    .io_read_bits_way_en(meta_io_read_bits_way_en),
    .io_write_ready(meta_io_write_ready),
    .io_write_valid(meta_io_write_valid),
    .io_write_bits_idx(meta_io_write_bits_idx),
    .io_write_bits_way_en(meta_io_write_bits_way_en),
    .io_write_bits_data_tag(meta_io_write_bits_data_tag),
    .io_write_bits_data_coh_state(meta_io_write_bits_data_coh_state),
    .io_resp_0_tag(meta_io_resp_0_tag),
    .io_resp_0_coh_state(meta_io_resp_0_coh_state)
  );
  Arbiter metaReadArb (
    .clk(metaReadArb_clk),
    .reset(metaReadArb_reset),
    .io_in_0_ready(metaReadArb_io_in_0_ready),
    .io_in_0_valid(metaReadArb_io_in_0_valid),
    .io_in_0_bits_idx(metaReadArb_io_in_0_bits_idx),
    .io_in_0_bits_way_en(metaReadArb_io_in_0_bits_way_en),
    .io_in_1_ready(metaReadArb_io_in_1_ready),
    .io_in_1_valid(metaReadArb_io_in_1_valid),
    .io_in_1_bits_idx(metaReadArb_io_in_1_bits_idx),
    .io_in_1_bits_way_en(metaReadArb_io_in_1_bits_way_en),
    .io_in_2_ready(metaReadArb_io_in_2_ready),
    .io_in_2_valid(metaReadArb_io_in_2_valid),
    .io_in_2_bits_idx(metaReadArb_io_in_2_bits_idx),
    .io_in_2_bits_way_en(metaReadArb_io_in_2_bits_way_en),
    .io_out_ready(metaReadArb_io_out_ready),
    .io_out_valid(metaReadArb_io_out_valid),
    .io_out_bits_idx(metaReadArb_io_out_bits_idx),
    .io_out_bits_way_en(metaReadArb_io_out_bits_way_en),
    .io_chosen(metaReadArb_io_chosen)
  );
  Arbiter_1 metaWriteArb (
    .clk(metaWriteArb_clk),
    .reset(metaWriteArb_reset),
    .io_in_0_ready(metaWriteArb_io_in_0_ready),
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_idx(metaWriteArb_io_in_0_bits_idx),
    .io_in_0_bits_way_en(metaWriteArb_io_in_0_bits_way_en),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_data_coh_state(metaWriteArb_io_in_0_bits_data_coh_state),
    .io_in_1_ready(metaWriteArb_io_in_1_ready),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_idx(metaWriteArb_io_in_1_bits_idx),
    .io_in_1_bits_way_en(metaWriteArb_io_in_1_bits_way_en),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_coh_state(metaWriteArb_io_in_1_bits_data_coh_state),
    .io_in_2_ready(metaWriteArb_io_in_2_ready),
    .io_in_2_valid(metaWriteArb_io_in_2_valid),
    .io_in_2_bits_idx(metaWriteArb_io_in_2_bits_idx),
    .io_in_2_bits_way_en(metaWriteArb_io_in_2_bits_way_en),
    .io_in_2_bits_data_tag(metaWriteArb_io_in_2_bits_data_tag),
    .io_in_2_bits_data_coh_state(metaWriteArb_io_in_2_bits_data_coh_state),
    .io_out_ready(metaWriteArb_io_out_ready),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_idx(metaWriteArb_io_out_bits_idx),
    .io_out_bits_way_en(metaWriteArb_io_out_bits_way_en),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_coh_state(metaWriteArb_io_out_bits_data_coh_state),
    .io_chosen(metaWriteArb_io_chosen)
  );
  DCacheDataArray data (
    .clk(data_clk),
    .reset(data_reset),
    .io_req_valid(data_io_req_valid),
    .io_req_bits_addr(data_io_req_bits_addr),
    .io_req_bits_write(data_io_req_bits_write),
    .io_req_bits_wdata(data_io_req_bits_wdata),
    .io_req_bits_wmask(data_io_req_bits_wmask),
    .io_req_bits_way_en(data_io_req_bits_way_en),
    .io_resp_0(data_io_resp_0)
  );
  Arbiter_2 dataArb (
    .clk(dataArb_clk),
    .reset(dataArb_reset),
    .io_in_0_ready(dataArb_io_in_0_ready),
    .io_in_0_valid(dataArb_io_in_0_valid),
    .io_in_0_bits_addr(dataArb_io_in_0_bits_addr),
    .io_in_0_bits_write(dataArb_io_in_0_bits_write),
    .io_in_0_bits_wdata(dataArb_io_in_0_bits_wdata),
    .io_in_0_bits_wmask(dataArb_io_in_0_bits_wmask),
    .io_in_0_bits_way_en(dataArb_io_in_0_bits_way_en),
    .io_in_1_ready(dataArb_io_in_1_ready),
    .io_in_1_valid(dataArb_io_in_1_valid),
    .io_in_1_bits_addr(dataArb_io_in_1_bits_addr),
    .io_in_1_bits_write(dataArb_io_in_1_bits_write),
    .io_in_1_bits_wdata(dataArb_io_in_1_bits_wdata),
    .io_in_1_bits_wmask(dataArb_io_in_1_bits_wmask),
    .io_in_1_bits_way_en(dataArb_io_in_1_bits_way_en),
    .io_in_2_ready(dataArb_io_in_2_ready),
    .io_in_2_valid(dataArb_io_in_2_valid),
    .io_in_2_bits_addr(dataArb_io_in_2_bits_addr),
    .io_in_2_bits_write(dataArb_io_in_2_bits_write),
    .io_in_2_bits_wdata(dataArb_io_in_2_bits_wdata),
    .io_in_2_bits_wmask(dataArb_io_in_2_bits_wmask),
    .io_in_2_bits_way_en(dataArb_io_in_2_bits_way_en),
    .io_in_3_ready(dataArb_io_in_3_ready),
    .io_in_3_valid(dataArb_io_in_3_valid),
    .io_in_3_bits_addr(dataArb_io_in_3_bits_addr),
    .io_in_3_bits_write(dataArb_io_in_3_bits_write),
    .io_in_3_bits_wdata(dataArb_io_in_3_bits_wdata),
    .io_in_3_bits_wmask(dataArb_io_in_3_bits_wmask),
    .io_in_3_bits_way_en(dataArb_io_in_3_bits_way_en),
    .io_out_ready(dataArb_io_out_ready),
    .io_out_valid(dataArb_io_out_valid),
    .io_out_bits_addr(dataArb_io_out_bits_addr),
    .io_out_bits_write(dataArb_io_out_bits_write),
    .io_out_bits_wdata(dataArb_io_out_bits_wdata),
    .io_out_bits_wmask(dataArb_io_out_bits_wmask),
    .io_out_bits_way_en(dataArb_io_out_bits_way_en),
    .io_chosen(dataArb_io_chosen)
  );
  TLB tlb (
    .clk(tlb_clk),
    .reset(tlb_reset),
    .io_req_ready(tlb_io_req_ready),
    .io_req_valid(tlb_io_req_valid),
    .io_req_bits_vpn(tlb_io_req_bits_vpn),
    .io_req_bits_passthrough(tlb_io_req_bits_passthrough),
    .io_req_bits_instruction(tlb_io_req_bits_instruction),
    .io_req_bits_store(tlb_io_req_bits_store),
    .io_resp_miss(tlb_io_resp_miss),
    .io_resp_ppn(tlb_io_resp_ppn),
    .io_resp_xcpt_ld(tlb_io_resp_xcpt_ld),
    .io_resp_xcpt_st(tlb_io_resp_xcpt_st),
    .io_resp_xcpt_if(tlb_io_resp_xcpt_if),
    .io_resp_cacheable(tlb_io_resp_cacheable),
    .io_ptw_req_ready(tlb_io_ptw_req_ready),
    .io_ptw_req_valid(tlb_io_ptw_req_valid),
    .io_ptw_req_bits_prv(tlb_io_ptw_req_bits_prv),
    .io_ptw_req_bits_pum(tlb_io_ptw_req_bits_pum),
    .io_ptw_req_bits_mxr(tlb_io_ptw_req_bits_mxr),
    .io_ptw_req_bits_addr(tlb_io_ptw_req_bits_addr),
    .io_ptw_req_bits_store(tlb_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(tlb_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(tlb_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_reserved_for_hardware(tlb_io_ptw_resp_bits_pte_reserved_for_hardware),
    .io_ptw_resp_bits_pte_ppn(tlb_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(tlb_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(tlb_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(tlb_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(tlb_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(tlb_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(tlb_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(tlb_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(tlb_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(tlb_io_ptw_resp_bits_pte_v),
    .io_ptw_ptbr_asid(tlb_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(tlb_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(tlb_io_ptw_invalidate),
    .io_ptw_status_debug(tlb_io_ptw_status_debug),
    .io_ptw_status_prv(tlb_io_ptw_status_prv),
    .io_ptw_status_sd(tlb_io_ptw_status_sd),
    .io_ptw_status_zero3(tlb_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(tlb_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(tlb_io_ptw_status_zero2),
    .io_ptw_status_vm(tlb_io_ptw_status_vm),
    .io_ptw_status_zero1(tlb_io_ptw_status_zero1),
    .io_ptw_status_mxr(tlb_io_ptw_status_mxr),
    .io_ptw_status_pum(tlb_io_ptw_status_pum),
    .io_ptw_status_mprv(tlb_io_ptw_status_mprv),
    .io_ptw_status_xs(tlb_io_ptw_status_xs),
    .io_ptw_status_fs(tlb_io_ptw_status_fs),
    .io_ptw_status_mpp(tlb_io_ptw_status_mpp),
    .io_ptw_status_hpp(tlb_io_ptw_status_hpp),
    .io_ptw_status_spp(tlb_io_ptw_status_spp),
    .io_ptw_status_mpie(tlb_io_ptw_status_mpie),
    .io_ptw_status_hpie(tlb_io_ptw_status_hpie),
    .io_ptw_status_spie(tlb_io_ptw_status_spie),
    .io_ptw_status_upie(tlb_io_ptw_status_upie),
    .io_ptw_status_mie(tlb_io_ptw_status_mie),
    .io_ptw_status_hie(tlb_io_ptw_status_hie),
    .io_ptw_status_sie(tlb_io_ptw_status_sie),
    .io_ptw_status_uie(tlb_io_ptw_status_uie)
  );
  assign io_cpu_req_ready = GEN_13;
  assign io_cpu_s2_nack = GEN_113;
  assign io_cpu_resp_valid = GEN_109;
  assign io_cpu_resp_bits_addr = s2_req_addr;
  assign io_cpu_resp_bits_tag = s2_req_tag;
  assign io_cpu_resp_bits_cmd = s2_req_cmd;
  assign io_cpu_resp_bits_typ = s2_req_typ;
  assign io_cpu_resp_bits_data = T_4496;
  assign io_cpu_resp_bits_replay = doUncachedResp;
  assign io_cpu_resp_bits_has_data = s2_read;
  assign io_cpu_resp_bits_data_word_bypass = s2_data_word[31:0];
  assign io_cpu_resp_bits_store_data = pstore1_data;
  assign io_cpu_replay_next = T_4443;
  assign io_cpu_xcpt_ma_ld = T_2903;
  assign io_cpu_xcpt_ma_st = T_2904;
  assign io_cpu_xcpt_pf_ld = T_2905;
  assign io_cpu_xcpt_pf_st = T_2906;
  assign io_cpu_ordered = T_4442;
  assign io_ptw_req_valid = tlb_io_ptw_req_valid;
  assign io_ptw_req_bits_prv = tlb_io_ptw_req_bits_prv;
  assign io_ptw_req_bits_pum = tlb_io_ptw_req_bits_pum;
  assign io_ptw_req_bits_mxr = tlb_io_ptw_req_bits_mxr;
  assign io_ptw_req_bits_addr = tlb_io_ptw_req_bits_addr;
  assign io_ptw_req_bits_store = tlb_io_ptw_req_bits_store;
  assign io_ptw_req_bits_fetch = tlb_io_ptw_req_bits_fetch;
  assign io_mem_acquire_valid = T_3731;
  assign io_mem_acquire_bits_addr_block = GEN_61;
  assign io_mem_acquire_bits_client_xact_id = GEN_62;
  assign io_mem_acquire_bits_addr_beat = GEN_63;
  assign io_mem_acquire_bits_is_builtin_type = GEN_64;
  assign io_mem_acquire_bits_a_type = GEN_65;
  assign io_mem_acquire_bits_union = GEN_66;
  assign io_mem_acquire_bits_data = GEN_67;
  assign io_mem_probe_ready = T_3932;
  assign io_mem_release_valid = GEN_86;
  assign io_mem_release_bits_addr_beat = writebackCount;
  assign io_mem_release_bits_addr_block = probe_bits_addr_block;
  assign io_mem_release_bits_client_xact_id = GEN_99;
  assign io_mem_release_bits_voluntary = GEN_100;
  assign io_mem_release_bits_r_type = GEN_101;
  assign io_mem_release_bits_data = s2_data;
  assign io_mem_grant_ready = 1'h1;
  assign io_mem_finish_valid = fq_io_deq_valid;
  assign io_mem_finish_bits_manager_xact_id = fq_io_deq_bits_manager_xact_id;
  assign io_mem_finish_bits_manager_id = fq_io_deq_bits_manager_id;
  assign fq_clk = clk;
  assign fq_reset = reset;
  assign fq_io_enq_valid = T_3867;
  assign fq_io_enq_bits_manager_xact_id = T_3891_manager_xact_id;
  assign fq_io_enq_bits_manager_id = T_3891_manager_id;
  assign fq_io_deq_ready = io_mem_finish_ready;
  assign T_1924 = refillDone;
  assign T_1928 = T_1927[0];
  assign T_1929 = T_1927[2];
  assign T_1930 = T_1928 ^ T_1929;
  assign T_1931 = T_1927[3];
  assign T_1932 = T_1930 ^ T_1931;
  assign T_1933 = T_1927[5];
  assign T_1934 = T_1932 ^ T_1933;
  assign T_1935 = T_1927[15:1];
  assign T_1936 = {T_1934,T_1935};
  assign GEN_2 = T_1924 ? T_1936 : T_1927;
  assign meta_clk = clk;
  assign meta_reset = reset;
  assign meta_io_read_valid = metaReadArb_io_out_valid;
  assign meta_io_read_bits_idx = metaReadArb_io_out_bits_idx;
  assign meta_io_read_bits_way_en = metaReadArb_io_out_bits_way_en;
  assign meta_io_write_valid = metaWriteArb_io_out_valid;
  assign meta_io_write_bits_idx = metaWriteArb_io_out_bits_idx;
  assign meta_io_write_bits_way_en = metaWriteArb_io_out_bits_way_en;
  assign meta_io_write_bits_data_tag = metaWriteArb_io_out_bits_data_tag;
  assign meta_io_write_bits_data_coh_state = metaWriteArb_io_out_bits_data_coh_state;
  assign metaReadArb_clk = clk;
  assign metaReadArb_reset = reset;
  assign metaReadArb_io_in_0_valid = flushing;
  assign metaReadArb_io_in_0_bits_idx = T_4508;
  assign metaReadArb_io_in_0_bits_way_en = 1'h1;
  assign metaReadArb_io_in_1_valid = T_3922;
  assign metaReadArb_io_in_1_bits_idx = io_mem_probe_bits_addr_block[6:0];
  assign metaReadArb_io_in_1_bits_way_en = 1'h1;
  assign metaReadArb_io_in_2_valid = io_cpu_req_valid;
  assign metaReadArb_io_in_2_bits_idx = T_2376;
  assign metaReadArb_io_in_2_bits_way_en = 1'h1;
  assign metaReadArb_io_out_ready = meta_io_read_ready;
  assign metaWriteArb_clk = clk;
  assign metaWriteArb_reset = reset;
  assign metaWriteArb_io_in_0_valid = T_3142;
  assign metaWriteArb_io_in_0_bits_idx = T_3143;
  assign metaWriteArb_io_in_0_bits_way_en = s2_victim_way[0];
  assign metaWriteArb_io_in_0_bits_data_tag = T_3211;
  assign metaWriteArb_io_in_0_bits_data_coh_state = T_3189_state;
  assign metaWriteArb_io_in_1_valid = refillDone;
  assign metaWriteArb_io_in_1_bits_idx = T_3143;
  assign metaWriteArb_io_in_1_bits_way_en = s2_victim_way[0];
  assign metaWriteArb_io_in_1_bits_data_tag = T_3211;
  assign metaWriteArb_io_in_1_bits_data_coh_state = T_3830_state;
  assign metaWriteArb_io_in_2_valid = T_4428;
  assign metaWriteArb_io_in_2_bits_idx = T_4432;
  assign metaWriteArb_io_in_2_bits_way_en = releaseWay[0];
  assign metaWriteArb_io_in_2_bits_data_tag = T_4436;
  assign metaWriteArb_io_in_2_bits_data_coh_state = newCoh_state;
  assign metaWriteArb_io_out_ready = meta_io_write_ready;
  assign data_clk = clk;
  assign data_reset = reset;
  assign data_io_req_valid = dataArb_io_out_valid;
  assign data_io_req_bits_addr = dataArb_io_out_bits_addr;
  assign data_io_req_bits_write = dataArb_io_out_bits_write;
  assign data_io_req_bits_wdata = dataArb_io_out_bits_wdata;
  assign data_io_req_bits_wmask = dataArb_io_out_bits_wmask;
  assign data_io_req_bits_way_en = dataArb_io_out_bits_way_en;
  assign dataArb_clk = clk;
  assign dataArb_reset = reset;
  assign dataArb_io_in_0_valid = T_2986;
  assign dataArb_io_in_0_bits_addr = T_3040[12:0];
  assign dataArb_io_in_0_bits_write = 1'h1;
  assign dataArb_io_in_0_bits_wdata = T_3043;
  assign dataArb_io_in_0_bits_wmask = T_3074[7:0];
  assign dataArb_io_in_0_bits_way_en = T_3041;
  assign dataArb_io_in_1_valid = T_3778;
  assign dataArb_io_in_1_bits_addr = T_3789[12:0];
  assign dataArb_io_in_1_bits_write = 1'h1;
  assign dataArb_io_in_1_bits_wdata = io_mem_grant_bits_data;
  assign dataArb_io_in_1_bits_wmask = 8'hff;
  assign dataArb_io_in_1_bits_way_en = s2_victim_way[0];
  assign dataArb_io_in_2_valid = T_4419;
  assign dataArb_io_in_2_bits_addr = T_4423[12:0];
  assign dataArb_io_in_2_bits_write = 1'h0;
  assign dataArb_io_in_2_bits_wdata = GEN_14;
  assign dataArb_io_in_2_bits_wmask = GEN_33;
  assign dataArb_io_in_2_bits_way_en = 1'h1;
  assign dataArb_io_in_3_valid = T_2359;
  assign dataArb_io_in_3_bits_addr = io_cpu_req_bits_addr[12:0];
  assign dataArb_io_in_3_bits_write = 1'h0;
  assign dataArb_io_in_3_bits_wdata = GEN_34;
  assign dataArb_io_in_3_bits_wmask = GEN_47;
  assign dataArb_io_in_3_bits_way_en = 1'h1;
  assign dataArb_io_out_ready = 1'h1;
  assign T_2218 = io_cpu_req_ready & io_cpu_req_valid;
  assign T_2220 = io_mem_probe_ready & io_mem_probe_valid;
  assign GEN_3 = T_2220 ? io_mem_probe_bits_addr_block : probe_bits_addr_block;
  assign GEN_4 = T_2220 ? io_mem_probe_bits_p_type : probe_bits_p_type;
  assign s1_nack = GEN_107;
  assign T_2247 = io_cpu_s1_kill == 1'h0;
  assign s1_valid_masked = s1_valid & T_2247;
  assign T_2249 = s1_nack == 1'h0;
  assign s1_valid_not_nacked = s1_valid_masked & T_2249;
  assign T_2316 = io_cpu_req_bits_addr[31:13];
  assign T_2317 = io_cpu_req_bits_addr[5:0];
  assign T_2318 = {T_2316,metaReadArb_io_out_bits_idx};
  assign T_2319 = {T_2318,T_2317};
  assign GEN_5 = metaReadArb_io_out_valid ? T_2319 : s1_req_addr;
  assign GEN_6 = metaReadArb_io_out_valid ? io_cpu_req_bits_tag : s1_req_tag;
  assign GEN_7 = metaReadArb_io_out_valid ? io_cpu_req_bits_cmd : s1_req_cmd;
  assign GEN_8 = metaReadArb_io_out_valid ? io_cpu_req_bits_typ : s1_req_typ;
  assign GEN_9 = metaReadArb_io_out_valid ? io_cpu_req_bits_phys : s1_req_phys;
  assign GEN_10 = metaReadArb_io_out_valid ? io_cpu_req_bits_data : s1_req_data;
  assign T_2320 = s1_req_cmd == 5'h0;
  assign T_2321 = s1_req_cmd == 5'h6;
  assign T_2322 = T_2320 | T_2321;
  assign T_2323 = s1_req_cmd == 5'h7;
  assign T_2324 = T_2322 | T_2323;
  assign T_2325 = s1_req_cmd[3];
  assign T_2326 = s1_req_cmd == 5'h4;
  assign T_2327 = T_2325 | T_2326;
  assign s1_read = T_2324 | T_2327;
  assign T_2328 = s1_req_cmd == 5'h1;
  assign T_2330 = T_2328 | T_2323;
  assign s1_write = T_2330 | T_2327;
  assign s1_readwrite = s1_read | s1_write;
  assign pstore1_valid = T_3001;
  assign T_2340 = release_state == 3'h2;
  assign T_2341 = release_state == 3'h3;
  assign inWriteback = T_2340 | T_2341;
  assign releaseWay = GEN_104;
  assign T_2343 = release_state == 3'h0;
  assign T_2345 = grant_wait == 1'h0;
  assign T_2346 = T_2343 & T_2345;
  assign T_2349 = T_2346 & T_2249;
  assign T_2350 = io_cpu_req_bits_cmd == 5'h0;
  assign T_2351 = io_cpu_req_bits_cmd == 5'h6;
  assign T_2352 = T_2350 | T_2351;
  assign T_2353 = io_cpu_req_bits_cmd == 5'h7;
  assign T_2354 = T_2352 | T_2353;
  assign T_2355 = io_cpu_req_bits_cmd[3];
  assign T_2356 = io_cpu_req_bits_cmd == 5'h4;
  assign T_2357 = T_2355 | T_2356;
  assign T_2358 = T_2354 | T_2357;
  assign T_2359 = io_cpu_req_valid & T_2358;
  assign T_2364 = dataArb_io_in_3_ready == 1'h0;
  assign T_2374 = T_2364 & T_2358;
  assign GEN_11 = T_2374 ? 1'h0 : T_2349;
  assign T_2376 = io_cpu_req_bits_addr[12:6];
  assign T_2380 = metaReadArb_io_in_2_ready == 1'h0;
  assign GEN_12 = T_2380 ? 1'h0 : GEN_11;
  assign tlb_clk = clk;
  assign tlb_reset = reset;
  assign tlb_io_req_valid = T_2382;
  assign tlb_io_req_bits_vpn = T_2383;
  assign tlb_io_req_bits_passthrough = s1_req_phys;
  assign tlb_io_req_bits_instruction = 1'h0;
  assign tlb_io_req_bits_store = s1_write;
  assign tlb_io_ptw_req_ready = io_ptw_req_ready;
  assign tlb_io_ptw_resp_valid = io_ptw_resp_valid;
  assign tlb_io_ptw_resp_bits_pte_reserved_for_hardware = io_ptw_resp_bits_pte_reserved_for_hardware;
  assign tlb_io_ptw_resp_bits_pte_ppn = io_ptw_resp_bits_pte_ppn;
  assign tlb_io_ptw_resp_bits_pte_reserved_for_software = io_ptw_resp_bits_pte_reserved_for_software;
  assign tlb_io_ptw_resp_bits_pte_d = io_ptw_resp_bits_pte_d;
  assign tlb_io_ptw_resp_bits_pte_a = io_ptw_resp_bits_pte_a;
  assign tlb_io_ptw_resp_bits_pte_g = io_ptw_resp_bits_pte_g;
  assign tlb_io_ptw_resp_bits_pte_u = io_ptw_resp_bits_pte_u;
  assign tlb_io_ptw_resp_bits_pte_x = io_ptw_resp_bits_pte_x;
  assign tlb_io_ptw_resp_bits_pte_w = io_ptw_resp_bits_pte_w;
  assign tlb_io_ptw_resp_bits_pte_r = io_ptw_resp_bits_pte_r;
  assign tlb_io_ptw_resp_bits_pte_v = io_ptw_resp_bits_pte_v;
  assign tlb_io_ptw_ptbr_asid = io_ptw_ptbr_asid;
  assign tlb_io_ptw_ptbr_ppn = io_ptw_ptbr_ppn;
  assign tlb_io_ptw_invalidate = io_ptw_invalidate;
  assign tlb_io_ptw_status_debug = io_ptw_status_debug;
  assign tlb_io_ptw_status_prv = io_ptw_status_prv;
  assign tlb_io_ptw_status_sd = io_ptw_status_sd;
  assign tlb_io_ptw_status_zero3 = io_ptw_status_zero3;
  assign tlb_io_ptw_status_sd_rv32 = io_ptw_status_sd_rv32;
  assign tlb_io_ptw_status_zero2 = io_ptw_status_zero2;
  assign tlb_io_ptw_status_vm = io_ptw_status_vm;
  assign tlb_io_ptw_status_zero1 = io_ptw_status_zero1;
  assign tlb_io_ptw_status_mxr = io_ptw_status_mxr;
  assign tlb_io_ptw_status_pum = io_ptw_status_pum;
  assign tlb_io_ptw_status_mprv = io_ptw_status_mprv;
  assign tlb_io_ptw_status_xs = io_ptw_status_xs;
  assign tlb_io_ptw_status_fs = io_ptw_status_fs;
  assign tlb_io_ptw_status_mpp = io_ptw_status_mpp;
  assign tlb_io_ptw_status_hpp = io_ptw_status_hpp;
  assign tlb_io_ptw_status_spp = io_ptw_status_spp;
  assign tlb_io_ptw_status_mpie = io_ptw_status_mpie;
  assign tlb_io_ptw_status_hpie = io_ptw_status_hpie;
  assign tlb_io_ptw_status_spie = io_ptw_status_spie;
  assign tlb_io_ptw_status_upie = io_ptw_status_upie;
  assign tlb_io_ptw_status_mie = io_ptw_status_mie;
  assign tlb_io_ptw_status_hie = io_ptw_status_hie;
  assign tlb_io_ptw_status_sie = io_ptw_status_sie;
  assign tlb_io_ptw_status_uie = io_ptw_status_uie;
  assign T_2382 = s1_valid_masked & s1_readwrite;
  assign T_2383 = s1_req_addr[31:12];
  assign T_2386 = tlb_io_req_ready == 1'h0;
  assign T_2388 = io_cpu_req_bits_phys == 1'h0;
  assign T_2389 = T_2386 & T_2388;
  assign GEN_13 = T_2389 ? 1'h0 : GEN_12;
  assign T_2391 = s1_valid & s1_readwrite;
  assign T_2392 = T_2391 & tlb_io_resp_miss;
  assign T_2394 = s1_req_addr[11:0];
  assign s1_paddr = {tlb_io_resp_ppn,T_2394};
  assign T_2395 = probe_bits_addr_block[25:7];
  assign T_2396 = s1_paddr[31:13];
  assign s1_tag = s1_probe ? T_2395 : T_2396;
  assign T_2397 = meta_io_resp_0_coh_state != 2'h0;
  assign T_2398 = meta_io_resp_0_tag == s1_tag;
  assign s1_hit_way = T_2397 & T_2398;
  assign T_2422_state = 2'h0;
  assign T_2446 = T_2398 ? meta_io_resp_0_coh_state : 2'h0;
  assign s1_hit_state_state = T_2446;
  assign s1_victim_way = 1'h0;
  assign T_2496 = s1_probe | s2_probe;
  assign T_2497 = release_state != 3'h0;
  assign releaseInFlight = T_2496 | T_2497;
  assign s2_valid_masked = s2_valid & T_2500;
  assign T_2568 = s1_valid_not_nacked | s1_flush_valid;
  assign T_2570 = tlb_io_resp_cacheable == 1'h0;
  assign GEN_15 = T_2568 ? s1_paddr : s2_req_addr;
  assign GEN_16 = T_2568 ? s1_req_tag : s2_req_tag;
  assign GEN_17 = T_2568 ? s1_req_cmd : s2_req_cmd;
  assign GEN_18 = T_2568 ? s1_req_typ : s2_req_typ;
  assign GEN_19 = T_2568 ? s1_req_phys : s2_req_phys;
  assign GEN_20 = T_2568 ? s1_req_data : s2_req_data;
  assign GEN_21 = T_2568 ? T_2570 : s2_uncached;
  assign T_2571 = s2_req_cmd == 5'h0;
  assign T_2572 = s2_req_cmd == 5'h6;
  assign T_2573 = T_2571 | T_2572;
  assign T_2574 = s2_req_cmd == 5'h7;
  assign T_2575 = T_2573 | T_2574;
  assign T_2576 = s2_req_cmd[3];
  assign T_2577 = s2_req_cmd == 5'h4;
  assign T_2578 = T_2576 | T_2577;
  assign s2_read = T_2575 | T_2578;
  assign T_2579 = s2_req_cmd == 5'h1;
  assign T_2581 = T_2579 | T_2574;
  assign s2_write = T_2581 | T_2578;
  assign s2_readwrite = s2_read | s2_write;
  assign T_2585 = s1_valid | inWriteback;
  assign GEN_22 = T_2585 ? data_io_resp_0 : s2_data;
  assign GEN_23 = s1_probe ? s1_hit_way : s2_probe_way;
  assign GEN_24 = s1_probe ? s1_hit_state_state : s2_probe_state_state;
  assign GEN_25 = s1_valid_not_nacked ? s1_hit_way : s2_hit_way;
  assign GEN_26 = s1_valid_not_nacked ? s1_hit_state_state : s2_hit_state_state;
  assign T_2635 = s2_req_cmd == 5'h3;
  assign T_2636 = s2_write | T_2635;
  assign T_2638 = T_2636 | T_2572;
  assign T_2639 = s2_hit_state_state == 2'h1;
  assign T_2640 = s2_hit_state_state == 2'h2;
  assign T_2641 = T_2639 | T_2640;
  assign s2_hit = T_2638 ? T_2641 : T_2641;
  assign T_2645 = s2_valid_masked & s2_readwrite;
  assign s2_valid_hit = T_2645 & s2_hit;
  assign T_2648 = s2_hit == 1'h0;
  assign T_2649 = T_2645 & T_2648;
  assign T_2650 = pstore1_valid | pstore2_valid;
  assign T_2652 = T_2650 == 1'h0;
  assign T_2653 = T_2649 & T_2652;
  assign T_2655 = release_ack_wait == 1'h0;
  assign s2_valid_miss = T_2653 & T_2655;
  assign T_2657 = s2_uncached == 1'h0;
  assign s2_valid_cached_miss = s2_valid_miss & T_2657;
  assign s2_victimize = s2_valid_cached_miss | s2_flush_valid;
  assign s2_valid_uncached = s2_valid_miss & s2_uncached;
  assign T_2658 = s2_hit_state_state != 2'h0;
  assign T_2660 = s2_flush_valid == 1'h0;
  assign T_2661 = T_2658 & T_2660;
  assign GEN_27 = T_2568 ? s1_victim_way : T_2663;
  assign T_2665 = 2'h1 << T_2663;
  assign s2_victim_way = T_2661 ? {{1'd0}, s2_hit_way} : T_2665;
  assign GEN_0 = GEN_28;
  assign GEN_28 = meta_io_resp_0_tag;
  assign GEN_29 = T_2568 ? GEN_0 : s2_victim_tag;
  assign GEN_1 = GEN_30;
  assign GEN_30 = meta_io_resp_0_coh_state;
  assign GEN_31 = T_2568 ? GEN_1 : T_2839_state;
  assign s2_victim_state_state = T_2661 ? s2_hit_state_state : T_2839_state;
  assign s2_victim_dirty = s2_victim_state_state == 2'h2;
  assign T_2883 = s2_valid_hit == 1'h0;
  assign T_2884 = s2_valid & T_2883;
  assign T_2885 = s2_valid_uncached & io_mem_acquire_ready;
  assign T_2887 = T_2885 == 1'h0;
  assign T_2888 = T_2884 & T_2887;
  assign GEN_32 = T_2884 ? 1'h1 : T_2392;
  assign T_2894 = s1_req_typ[1:0];
  assign T_2896 = 4'h1 << T_2894;
  assign T_2898 = T_2896 - 4'h1;
  assign T_2899 = T_2898[3:0];
  assign T_2900 = T_2899[1:0];
  assign GEN_123 = {{30'd0}, T_2900};
  assign T_2901 = s1_req_addr & GEN_123;
  assign misaligned = T_2901 != 32'h0;
  assign T_2903 = s1_read & misaligned;
  assign T_2904 = s1_write & misaligned;
  assign T_2905 = s1_read & tlb_io_resp_xcpt_ld;
  assign T_2906 = s1_write & tlb_io_resp_xcpt_st;
  assign T_2907 = io_cpu_xcpt_ma_ld | io_cpu_xcpt_ma_st;
  assign T_2908 = T_2907 | io_cpu_xcpt_pf_ld;
  assign T_2909 = T_2908 | io_cpu_xcpt_pf_st;
  assign T_2911 = T_2910 & s2_valid_masked;
  assign T_2913 = T_2911 == 1'h0;
  assign T_2914 = T_2913 | reset;
  assign T_2916 = T_2914 == 1'h0;
  assign lrscValid = lrscCount > 5'h0;
  assign T_2933 = lrscCount - 5'h1;
  assign T_2934 = T_2933[4:0];
  assign GEN_35 = lrscValid ? T_2934 : lrscCount;
  assign GEN_36 = io_cpu_invalidate_lr ? 5'h0 : GEN_35;
  assign T_2938 = s1_valid_not_nacked & s1_write;
  assign GEN_37 = T_2938 ? s1_req_cmd : pstore1_cmd;
  assign GEN_38 = T_2938 ? s1_req_typ : pstore1_typ;
  assign GEN_39 = T_2938 ? s1_paddr : pstore1_addr;
  assign GEN_40 = T_2938 ? io_cpu_s1_data : pstore1_data;
  assign GEN_41 = T_2938 ? s1_hit_way : pstore1_way;
  assign T_2943 = pstore1_typ[1:0];
  assign T_2945 = T_2943 == 2'h0;
  assign T_2946 = pstore1_data[7:0];
  assign T_2947 = {T_2946,T_2946};
  assign T_2948 = {T_2947,T_2947};
  assign T_2950 = T_2943 == 2'h1;
  assign T_2951 = pstore1_data[15:0];
  assign T_2952 = {T_2951,T_2951};
  assign T_2953 = T_2950 ? T_2952 : pstore1_data;
  assign T_2954 = T_2945 ? T_2948 : T_2953;
  assign pstore1_storegen_data = T_2954;
  assign pstore_drain_opportunistic = T_2359 == 1'h0;
  assign pstore_drain_on_miss = releaseInFlight | io_cpu_s2_nack;
  assign T_2985 = pstore_drain_opportunistic | pstore_drain_on_miss;
  assign T_2986 = T_2650 & T_2985;
  assign T_2987 = s2_valid_hit & s2_write;
  assign T_2994 = T_2987 == 1'h0;
  assign T_2996 = T_2992 == 1'h0;
  assign T_2997 = T_2994 | T_2996;
  assign T_2998 = T_2997 | reset;
  assign T_3000 = T_2998 == 1'h0;
  assign T_3001 = T_2987 | T_2992;
  assign T_3002 = T_3001 & pstore2_valid;
  assign T_3004 = T_2986 == 1'h0;
  assign T_3005 = T_3002 & T_3004;
  assign T_3007 = pstore2_valid == T_2986;
  assign advance_pstore1 = pstore1_valid & T_3007;
  assign T_3010 = pstore2_valid & T_3004;
  assign T_3011 = T_3010 | advance_pstore1;
  assign GEN_42 = advance_pstore1 ? pstore1_addr : pstore2_addr;
  assign GEN_43 = advance_pstore1 ? pstore1_way : pstore2_way;
  assign GEN_44 = advance_pstore1 ? pstore1_storegen_data : pstore2_storegen_data;
  assign T_3013 = pstore1_addr[0];
  assign T_3017 = T_2943 >= 2'h1;
  assign T_3021 = T_3013 | T_3017;
  assign T_3024 = T_3013 ? 1'h0 : 1'h1;
  assign T_3025 = {T_3021,T_3024};
  assign T_3026 = pstore1_addr[1];
  assign T_3028 = T_3026 ? T_3025 : 2'h0;
  assign T_3030 = T_2943 >= 2'h2;
  assign T_3033 = T_3030 ? 2'h3 : 2'h0;
  assign T_3034 = T_3028 | T_3033;
  assign T_3037 = T_3026 ? 2'h0 : T_3025;
  assign T_3038 = {T_3034,T_3037};
  assign GEN_45 = advance_pstore1 ? T_3038 : pstore2_storegen_mask;
  assign T_3040 = pstore2_valid ? pstore2_addr : pstore1_addr;
  assign T_3041 = pstore2_valid ? pstore2_way : pstore1_way;
  assign T_3042 = pstore2_valid ? pstore2_storegen_data : pstore1_storegen_data;
  assign T_3043 = {T_3042,T_3042};
  assign T_3045 = T_3040[2];
  assign GEN_124 = {{2'd0}, T_3045};
  assign pstore_mask_shift = GEN_124 << 2;
  assign T_3073 = pstore2_valid ? pstore2_storegen_mask : T_3038;
  assign GEN_125 = {{7'd0}, T_3073};
  assign T_3074 = GEN_125 << pstore_mask_shift;
  assign s1_idx = s1_req_addr[12:2];
  assign T_3075 = pstore1_addr[12:2];
  assign T_3076 = T_3075 == s1_idx;
  assign T_3077 = pstore1_valid & T_3076;
  assign T_3078 = pstore2_addr[12:2];
  assign T_3079 = T_3078 == s1_idx;
  assign T_3080 = pstore2_valid & T_3079;
  assign T_3081 = T_3077 | T_3080;
  assign s1_raw_hazard = s1_read & T_3081;
  assign T_3082 = s1_valid & s1_raw_hazard;
  assign GEN_46 = T_3082 ? 1'h1 : GEN_32;
  assign T_3091 = s2_write ? 2'h2 : s2_hit_state_state;
  assign s2_new_hit_state_state = T_3091;
  assign T_3135 = s2_hit_state_state == s2_new_hit_state_state;
  assign T_3137 = T_3135 == 1'h0;
  assign T_3138 = s2_valid_hit & T_3137;
  assign T_3140 = s2_victim_dirty == 1'h0;
  assign T_3141 = s2_victimize & T_3140;
  assign T_3142 = T_3138 | T_3141;
  assign T_3143 = s2_req_addr[12:6];
  assign T_3167_state = 2'h0;
  assign T_3189_state = s2_hit ? s2_new_hit_state_state : T_3167_state;
  assign T_3211 = s2_req_addr[31:13];
  assign T_3213 = s2_req_addr[31:6];
  assign T_3228 = {s2_req_cmd,1'h1};
  assign cachedGetMessage_addr_block = T_3213;
  assign cachedGetMessage_client_xact_id = 1'h0;
  assign cachedGetMessage_addr_beat = 3'h0;
  assign cachedGetMessage_is_builtin_type = 1'h0;
  assign cachedGetMessage_a_type = {{2'd0}, T_2638};
  assign cachedGetMessage_union = {{6'd0}, T_3228};
  assign cachedGetMessage_data = 64'h0;
  assign T_3288 = s2_req_addr[5:3];
  assign T_3289 = s2_req_addr[2:0];
  assign T_3330 = {T_3289,s2_req_typ};
  assign T_3331 = {T_3330,6'h0};
  assign uncachedGetMessage_addr_block = T_3213;
  assign uncachedGetMessage_client_xact_id = 1'h0;
  assign uncachedGetMessage_addr_beat = T_3288;
  assign uncachedGetMessage_is_builtin_type = 1'h1;
  assign uncachedGetMessage_a_type = 3'h0;
  assign uncachedGetMessage_union = T_3331;
  assign uncachedGetMessage_data = 64'h0;
  assign uncachedPutOffset = s2_req_addr[2];
  assign T_3430 = {T_2954,T_2954};
  assign GEN_126 = {{2'd0}, uncachedPutOffset};
  assign T_3458 = GEN_126 << 2;
  assign GEN_127 = {{7'd0}, T_3038};
  assign T_3459 = GEN_127 << T_3458;
  assign T_3496 = T_3459[7:0];
  assign T_3506 = {T_3496,1'h0};
  assign T_3526 = {{3'd0}, T_3506};
  assign uncachedPutMessage_addr_block = T_3213;
  assign uncachedPutMessage_client_xact_id = 1'h0;
  assign uncachedPutMessage_addr_beat = T_3288;
  assign uncachedPutMessage_is_builtin_type = 1'h1;
  assign uncachedPutMessage_a_type = 3'h2;
  assign uncachedPutMessage_union = T_3526;
  assign uncachedPutMessage_data = T_3430;
  assign T_3642 = {T_3330,T_3228};
  assign uncachedPutAtomicMessage_addr_block = T_3213;
  assign uncachedPutAtomicMessage_client_xact_id = 1'h0;
  assign uncachedPutAtomicMessage_addr_beat = T_3288;
  assign uncachedPutAtomicMessage_is_builtin_type = 1'h1;
  assign uncachedPutAtomicMessage_a_type = 3'h4;
  assign uncachedPutAtomicMessage_union = T_3642;
  assign uncachedPutAtomicMessage_data = T_3430;
  assign T_3729 = s2_valid_cached_miss & T_3140;
  assign T_3730 = T_3729 | s2_valid_uncached;
  assign T_3731 = T_3730 & fq_io_enq_ready;
  assign T_3733 = s2_valid_masked == 1'h0;
  assign T_3736 = T_2658 == 1'h0;
  assign T_3737 = T_3733 | T_3736;
  assign T_3738 = T_3737 | reset;
  assign T_3740 = T_3738 == 1'h0;
  assign GEN_54 = s2_write ? uncachedPutMessage_addr_block : uncachedGetMessage_addr_block;
  assign GEN_55 = s2_write ? uncachedPutMessage_client_xact_id : uncachedGetMessage_client_xact_id;
  assign GEN_56 = s2_write ? uncachedPutMessage_addr_beat : uncachedGetMessage_addr_beat;
  assign GEN_57 = s2_write ? uncachedPutMessage_is_builtin_type : uncachedGetMessage_is_builtin_type;
  assign GEN_58 = s2_write ? uncachedPutMessage_a_type : uncachedGetMessage_a_type;
  assign GEN_59 = s2_write ? uncachedPutMessage_union : uncachedGetMessage_union;
  assign GEN_60 = s2_write ? uncachedPutMessage_data : uncachedGetMessage_data;
  assign GEN_61 = s2_uncached ? GEN_54 : cachedGetMessage_addr_block;
  assign GEN_62 = s2_uncached ? GEN_55 : cachedGetMessage_client_xact_id;
  assign GEN_63 = s2_uncached ? GEN_56 : cachedGetMessage_addr_beat;
  assign GEN_64 = s2_uncached ? GEN_57 : cachedGetMessage_is_builtin_type;
  assign GEN_65 = s2_uncached ? GEN_58 : cachedGetMessage_a_type;
  assign GEN_66 = s2_uncached ? GEN_59 : cachedGetMessage_union;
  assign GEN_67 = s2_uncached ? GEN_60 : cachedGetMessage_data;
  assign T_3741 = io_mem_acquire_ready & io_mem_acquire_valid;
  assign GEN_68 = T_3741 ? 1'h1 : grant_wait;
  assign T_3750_0 = 3'h5;
  assign GEN_128 = {{1'd0}, T_3750_0};
  assign T_3752 = io_mem_grant_bits_g_type == GEN_128;
  assign T_3753 = io_mem_grant_bits_g_type == 4'h0;
  assign T_3754 = io_mem_grant_bits_is_builtin_type ? T_3752 : T_3753;
  assign grantIsVoluntary = io_mem_grant_bits_is_builtin_type & T_3753;
  assign T_3758 = T_3754 == 1'h0;
  assign T_3760 = grantIsVoluntary == 1'h0;
  assign grantIsUncached = T_3758 & T_3760;
  assign T_3761 = grantIsVoluntary & release_ack_wait;
  assign T_3762 = grant_wait | T_3761;
  assign T_3763 = T_3762 | reset;
  assign T_3765 = T_3763 == 1'h0;
  assign GEN_69 = grantIsUncached ? io_mem_grant_bits_data : GEN_22;
  assign GEN_70 = grantIsVoluntary ? 1'h0 : release_ack_wait;
  assign GEN_71 = io_mem_grant_valid ? GEN_69 : GEN_22;
  assign GEN_72 = io_mem_grant_valid ? GEN_70 : release_ack_wait;
  assign T_3767 = io_mem_grant_ready & io_mem_grant_valid;
  assign T_3768 = T_3767 & T_3754;
  assign T_3771 = refillCount == 3'h7;
  assign T_3773 = refillCount + 3'h1;
  assign T_3774 = T_3773[2:0];
  assign GEN_73 = T_3768 ? T_3774 : refillCount;
  assign refillDone = T_3768 & T_3771;
  assign grantDone = refillDone | grantIsUncached;
  assign T_3776 = T_3767 & grantDone;
  assign GEN_74 = T_3776 ? 1'h0 : GEN_68;
  assign T_3778 = T_3754 & io_mem_grant_valid;
  assign T_3781 = dataArb_io_in_1_valid == 1'h0;
  assign T_3782 = dataArb_io_in_1_ready | T_3781;
  assign T_3783 = T_3782 | reset;
  assign T_3785 = T_3783 == 1'h0;
  assign T_3788 = {T_3213,io_mem_grant_bits_addr_beat};
  assign GEN_129 = {{3'd0}, T_3788};
  assign T_3789 = GEN_129 << 3;
  assign T_3793 = metaWriteArb_io_in_1_valid == 1'h0;
  assign T_3794 = T_3793 | metaWriteArb_io_in_1_ready;
  assign T_3795 = T_3794 | reset;
  assign T_3797 = T_3795 == 1'h0;
  assign T_3806 = s2_write ? 2'h2 : 2'h1;
  assign T_3807 = io_mem_grant_bits_is_builtin_type ? 2'h0 : T_3806;
  assign T_3830_state = T_3807;
  assign T_3863 = T_3767 & T_3760;
  assign T_3866 = T_3758 | refillDone;
  assign T_3867 = T_3863 & T_3866;
  assign T_3891_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign T_3891_manager_id = io_mem_grant_bits_manager_id;
  assign T_3914 = fq_io_enq_ready | reset;
  assign T_3916 = T_3914 == 1'h0;
  assign T_3918 = releaseInFlight | lrscValid;
  assign T_3921 = T_3918 == 1'h0;
  assign T_3922 = io_mem_probe_valid & T_3921;
  assign T_3925 = metaReadArb_io_in_1_ready & T_3921;
  assign T_3927 = s1_valid == 1'h0;
  assign T_3928 = T_3925 & T_3927;
  assign T_3930 = s2_valid == 1'h0;
  assign T_3931 = T_3930 | s2_valid_hit;
  assign T_3932 = T_3928 & T_3931;
  assign T_3935 = io_mem_release_ready & io_mem_release_valid;
  assign T_3936 = T_3935 & inWriteback;
  assign T_3939 = writebackCount == 3'h7;
  assign T_3941 = writebackCount + 3'h1;
  assign T_3942 = T_3941[2:0];
  assign GEN_76 = T_3936 ? T_3942 : writebackCount;
  assign writebackDone = T_3936 & T_3939;
  assign T_3945 = inWriteback == 1'h0;
  assign T_3946 = T_3935 & T_3945;
  assign releaseDone = writebackDone | T_3946;
  assign T_3948 = io_mem_release_ready == 1'h0;
  assign releaseRejected = io_mem_release_valid & T_3948;
  assign T_3949 = dataArb_io_in_2_ready & dataArb_io_in_2_valid;
  assign T_3951 = releaseRejected == 1'h0;
  assign T_3952 = s1_release_data_valid & T_3951;
  assign T_3954 = {1'h0,writebackCount};
  assign T_3957 = {1'h0,s2_release_data_valid};
  assign GEN_130 = {{1'd0}, s1_release_data_valid};
  assign T_3958 = GEN_130 + T_3957;
  assign T_3959 = T_3958[1:0];
  assign T_3960 = releaseRejected ? 2'h0 : T_3959;
  assign GEN_131 = {{2'd0}, T_3960};
  assign T_3961 = T_3954 + GEN_131;
  assign releaseDataBeat = T_3961[3:0];
  assign T_3985_state = 2'h0;
  assign T_4010 = T_3985_state == 2'h2;
  assign T_4011 = T_4010 ? 3'h0 : 3'h3;
  assign T_4040 = 2'h2 == probe_bits_p_type;
  assign T_4041 = T_4040 ? T_4011 : 3'h3;
  assign T_4042 = 2'h1 == probe_bits_p_type;
  assign T_4043 = T_4042 ? T_4011 : T_4041;
  assign T_4044 = 2'h0 == probe_bits_p_type;
  assign T_4045 = T_4044 ? T_4011 : T_4043;
  assign T_4074_addr_beat = 3'h0;
  assign T_4074_addr_block = probe_bits_addr_block;
  assign T_4074_client_xact_id = 1'h0;
  assign T_4074_voluntary = 1'h0;
  assign T_4074_r_type = T_4045;
  assign T_4074_data = 64'h0;
  assign T_4107 = s2_victim_dirty ? 3'h0 : 3'h3;
  assign voluntaryReleaseMessage_addr_beat = 3'h0;
  assign voluntaryReleaseMessage_addr_block = 26'h0;
  assign voluntaryReleaseMessage_client_xact_id = 1'h0;
  assign voluntaryReleaseMessage_voluntary = 1'h1;
  assign voluntaryReleaseMessage_r_type = T_4107;
  assign voluntaryReleaseMessage_data = 64'h0;
  assign voluntaryNewCoh_state = 2'h0;
  assign T_4221 = s2_probe_state_state == 2'h2;
  assign T_4222 = T_4221 ? 3'h0 : 3'h3;
  assign T_4252 = T_4040 ? T_4222 : 3'h3;
  assign T_4254 = T_4042 ? T_4222 : T_4252;
  assign T_4256 = T_4044 ? T_4222 : T_4254;
  assign probeResponseMessage_addr_beat = 3'h0;
  assign probeResponseMessage_addr_block = probe_bits_addr_block;
  assign probeResponseMessage_client_xact_id = 1'h0;
  assign probeResponseMessage_voluntary = 1'h0;
  assign probeResponseMessage_r_type = T_4256;
  assign probeResponseMessage_data = 64'h0;
  assign T_4312 = T_4040 ? 2'h0 : s2_probe_state_state;
  assign T_4314 = T_4042 ? 2'h0 : T_4312;
  assign T_4316 = T_4044 ? 2'h0 : T_4314;
  assign probeNewCoh_state = T_4316;
  assign newCoh_state = GEN_103;
  assign T_4381 = s2_victimize & s2_victim_dirty;
  assign T_4385 = T_3736 | reset;
  assign T_4387 = T_4385 == 1'h0;
  assign T_4389 = {s2_victim_tag,T_3143};
  assign GEN_77 = T_4381 ? 3'h2 : release_state;
  assign GEN_78 = T_4381 ? T_4389 : GEN_3;
  assign GEN_79 = T_4221 ? 3'h3 : GEN_77;
  assign T_4391 = s2_probe_state_state != 2'h0;
  assign T_4393 = T_4221 == 1'h0;
  assign T_4394 = T_4393 & T_4391;
  assign GEN_80 = T_4394 ? 3'h4 : GEN_79;
  assign T_4398 = T_4391 == 1'h0;
  assign T_4399 = T_4393 & T_4398;
  assign GEN_81 = T_4399 ? 1'h1 : s2_release_data_valid;
  assign GEN_82 = T_4399 ? 3'h5 : GEN_80;
  assign GEN_83 = s2_probe ? GEN_82 : GEN_77;
  assign GEN_84 = s2_probe ? GEN_81 : s2_release_data_valid;
  assign GEN_85 = releaseDone ? 3'h0 : GEN_83;
  assign T_4401 = release_state == 3'h5;
  assign T_4402 = release_state == 3'h4;
  assign T_4403 = T_4401 | T_4402;
  assign GEN_86 = T_4403 ? 1'h1 : GEN_84;
  assign T_4407 = T_4402 | T_2341;
  assign GEN_87 = releaseDone ? 3'h7 : GEN_85;
  assign GEN_90 = T_4407 ? probeResponseMessage_client_xact_id : T_4074_client_xact_id;
  assign GEN_91 = T_4407 ? probeResponseMessage_voluntary : T_4074_voluntary;
  assign GEN_92 = T_4407 ? probeResponseMessage_r_type : T_4074_r_type;
  assign GEN_94 = T_4407 ? GEN_87 : GEN_85;
  assign T_4409 = release_state == 3'h6;
  assign T_4410 = T_2340 | T_4409;
  assign GEN_95 = releaseDone ? 3'h6 : GEN_94;
  assign GEN_96 = releaseDone ? 1'h1 : GEN_72;
  assign GEN_99 = T_4410 ? voluntaryReleaseMessage_client_xact_id : GEN_90;
  assign GEN_100 = T_4410 ? voluntaryReleaseMessage_voluntary : GEN_91;
  assign GEN_101 = T_4410 ? voluntaryReleaseMessage_r_type : GEN_92;
  assign GEN_103 = T_4410 ? voluntaryNewCoh_state : probeNewCoh_state;
  assign GEN_104 = T_4410 ? s2_victim_way : {{1'd0}, s2_probe_way};
  assign GEN_105 = T_4410 ? GEN_95 : GEN_94;
  assign GEN_106 = T_4410 ? GEN_96 : GEN_72;
  assign T_4414 = T_3935 == 1'h0;
  assign T_4415 = s2_probe & T_4414;
  assign GEN_107 = T_4415 ? 1'h1 : GEN_46;
  assign T_4418 = releaseDataBeat < 4'h8;
  assign T_4419 = inWriteback & T_4418;
  assign T_4421 = releaseDataBeat[2:0];
  assign T_4422 = {io_mem_release_bits_addr_block,T_4421};
  assign GEN_132 = {{3'd0}, T_4422};
  assign T_4423 = GEN_132 << 3;
  assign T_4427 = release_state == 3'h7;
  assign T_4428 = T_4409 | T_4427;
  assign T_4430 = {io_mem_release_bits_addr_block,io_mem_release_bits_addr_beat};
  assign T_4431 = {T_4430,3'h0};
  assign T_4432 = T_4431[12:6];
  assign T_4436 = T_4431[31:13];
  assign T_4437 = metaWriteArb_io_in_2_ready & metaWriteArb_io_in_2_valid;
  assign GEN_108 = T_4437 ? 3'h0 : GEN_105;
  assign T_4439 = s1_valid | s2_valid;
  assign T_4440 = T_4439 | grant_wait;
  assign T_4442 = T_4440 == 1'h0;
  assign T_4443 = io_mem_grant_valid & grantIsUncached;
  assign T_4446 = T_2883 | reset;
  assign T_4448 = T_4446 == 1'h0;
  assign GEN_109 = doUncachedResp ? 1'h1 : s2_valid_hit;
  assign T_4452 = {uncachedPutOffset,5'h0};
  assign s2_data_word = s2_data >> T_4452;
  assign T_4453 = s2_req_typ[1:0];
  assign T_4454 = $signed(s2_req_typ);
  assign T_4456 = $signed(T_4454) >= $signed(3'sh0);
  assign T_4457 = s2_req_addr[1];
  assign T_4458 = s2_data_word[31:16];
  assign T_4459 = s2_data_word[15:0];
  assign T_4460 = T_4457 ? T_4458 : T_4459;
  assign T_4466 = T_4453 == 2'h1;
  assign T_4468 = T_4460[15];
  assign T_4469 = T_4456 & T_4468;
  assign T_4473 = T_4469 ? 16'hffff : 16'h0;
  assign T_4475 = T_4466 ? T_4473 : T_4458;
  assign T_4476 = {T_4475,T_4460};
  assign T_4477 = s2_req_addr[0];
  assign T_4478 = T_4476[15:8];
  assign T_4479 = T_4476[7:0];
  assign T_4480 = T_4477 ? T_4478 : T_4479;
  assign T_4486 = T_4453 == 2'h0;
  assign T_4488 = T_4480[7];
  assign T_4489 = T_4456 & T_4488;
  assign T_4493 = T_4489 ? 24'hffffff : 24'h0;
  assign T_4494 = T_4476[31:8];
  assign T_4495 = T_4486 ? T_4493 : T_4494;
  assign T_4496 = {T_4495,T_4480};
  assign T_4498 = s1_valid_masked & s1_read;
  assign T_4499 = T_4498 & s1_write;
  assign T_4501 = T_4499 == 1'h0;
  assign T_4502 = T_4501 | reset;
  assign T_4504 = T_4502 == 1'h0;
  assign GEN_111 = T_3741 ? 1'h0 : flushed;
  assign T_4511 = s2_req_cmd == 5'h5;
  assign T_4512 = s2_valid_masked & T_4511;
  assign T_4514 = flushed == 1'h0;
  assign GEN_112 = T_4514 ? T_2655 : flushing;
  assign GEN_113 = T_4512 ? T_4514 : T_2888;
  assign GEN_114 = T_4512 ? GEN_112 : flushing;
  assign T_4519 = metaReadArb_io_in_0_ready & metaReadArb_io_in_0_valid;
  assign T_4521 = s1_flush_valid == 1'h0;
  assign T_4522 = T_4519 & T_4521;
  assign T_4525 = T_4522 & T_2660;
  assign T_4527 = T_4525 & T_2343;
  assign T_4530 = T_4527 & T_2655;
  assign T_4535 = T_4508 == 7'h7f;
  assign T_4537 = T_4508 + 7'h1;
  assign T_4538 = T_4537[6:0];
  assign GEN_115 = T_4535 ? 1'h1 : GEN_111;
  assign GEN_116 = s2_flush_valid ? T_4538 : T_4508;
  assign GEN_117 = s2_flush_valid ? GEN_115 : GEN_111;
  assign T_4541 = flushed & T_2343;
  assign T_4544 = T_4541 & T_2655;
  assign GEN_118 = T_4544 ? 1'h0 : GEN_114;
  assign GEN_120 = flushing ? GEN_116 : T_4508;
  assign GEN_121 = flushing ? GEN_117 : GEN_111;
  assign GEN_122 = flushing ? GEN_118 : GEN_114;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_48 = {1{$random}};
  T_1927 = GEN_48[15:0];
  `endif
  `ifdef RANDOMIZE
  GEN_49 = {1{$random}};
  s1_valid = GEN_49[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_50 = {1{$random}};
  s1_probe = GEN_50[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_51 = {1{$random}};
  probe_bits_addr_block = GEN_51[25:0];
  `endif
  `ifdef RANDOMIZE
  GEN_52 = {1{$random}};
  probe_bits_p_type = GEN_52[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_53 = {1{$random}};
  s1_req_addr = GEN_53[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_75 = {1{$random}};
  s1_req_tag = GEN_75[8:0];
  `endif
  `ifdef RANDOMIZE
  GEN_88 = {1{$random}};
  s1_req_cmd = GEN_88[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_89 = {1{$random}};
  s1_req_typ = GEN_89[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_93 = {1{$random}};
  s1_req_phys = GEN_93[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_97 = {1{$random}};
  s1_req_data = GEN_97[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_98 = {1{$random}};
  s1_flush_valid = GEN_98[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_102 = {1{$random}};
  grant_wait = GEN_102[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_110 = {1{$random}};
  release_ack_wait = GEN_110[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_119 = {1{$random}};
  release_state = GEN_119[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_133 = {1{$random}};
  pstore2_valid = GEN_133[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_134 = {1{$random}};
  s2_valid = GEN_134[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_135 = {1{$random}};
  s2_probe = GEN_135[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_136 = {1{$random}};
  T_2500 = GEN_136[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_137 = {1{$random}};
  s2_req_addr = GEN_137[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_138 = {1{$random}};
  s2_req_tag = GEN_138[8:0];
  `endif
  `ifdef RANDOMIZE
  GEN_139 = {1{$random}};
  s2_req_cmd = GEN_139[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_140 = {1{$random}};
  s2_req_typ = GEN_140[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_141 = {1{$random}};
  s2_req_phys = GEN_141[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_142 = {1{$random}};
  s2_req_data = GEN_142[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_143 = {1{$random}};
  s2_uncached = GEN_143[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_144 = {1{$random}};
  s2_flush_valid = GEN_144[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_145 = {2{$random}};
  s2_data = GEN_145[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_146 = {1{$random}};
  s2_probe_way = GEN_146[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_147 = {1{$random}};
  s2_probe_state_state = GEN_147[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_148 = {1{$random}};
  s2_hit_way = GEN_148[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_149 = {1{$random}};
  s2_hit_state_state = GEN_149[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_150 = {1{$random}};
  T_2663 = GEN_150[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_151 = {1{$random}};
  s2_victim_tag = GEN_151[18:0];
  `endif
  `ifdef RANDOMIZE
  GEN_152 = {1{$random}};
  T_2839_state = GEN_152[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_153 = {1{$random}};
  T_2910 = GEN_153[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_154 = {1{$random}};
  lrscCount = GEN_154[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_155 = {1{$random}};
  lrscAddr = GEN_155[25:0];
  `endif
  `ifdef RANDOMIZE
  GEN_156 = {1{$random}};
  pstore1_cmd = GEN_156[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_157 = {1{$random}};
  pstore1_typ = GEN_157[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_158 = {1{$random}};
  pstore1_addr = GEN_158[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_159 = {1{$random}};
  pstore1_data = GEN_159[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_160 = {1{$random}};
  pstore1_way = GEN_160[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_161 = {1{$random}};
  T_2992 = GEN_161[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_162 = {1{$random}};
  pstore2_addr = GEN_162[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_163 = {1{$random}};
  pstore2_way = GEN_163[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_164 = {1{$random}};
  pstore2_storegen_data = GEN_164[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_165 = {1{$random}};
  pstore2_storegen_mask = GEN_165[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_166 = {1{$random}};
  refillCount = GEN_166[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_167 = {1{$random}};
  writebackCount = GEN_167[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_168 = {1{$random}};
  s1_release_data_valid = GEN_168[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_169 = {1{$random}};
  s2_release_data_valid = GEN_169[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_170 = {1{$random}};
  doUncachedResp = GEN_170[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_171 = {1{$random}};
  flushed = GEN_171[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_172 = {1{$random}};
  flushing = GEN_172[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_173 = {1{$random}};
  T_4508 = GEN_173[6:0];
  `endif
  `ifdef RANDOMIZE
  GEN_174 = {2{$random}};
  GEN_14 = GEN_174[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_175 = {1{$random}};
  GEN_33 = GEN_175[7:0];
  `endif
  `ifdef RANDOMIZE
  GEN_176 = {2{$random}};
  GEN_34 = GEN_176[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_177 = {1{$random}};
  GEN_47 = GEN_177[7:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1927 <= 16'h1;
    end else begin
      if(T_1924) begin
        T_1927 <= T_1936;
      end
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T_2218;
    end
    if(reset) begin
      s1_probe <= 1'h0;
    end else begin
      s1_probe <= T_2220;
    end
    if(1'h0) begin
    end else begin
      if(T_4381) begin
        probe_bits_addr_block <= T_4389;
      end else begin
        if(T_2220) begin
          probe_bits_addr_block <= io_mem_probe_bits_addr_block;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2220) begin
        probe_bits_p_type <= io_mem_probe_bits_p_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(metaReadArb_io_out_valid) begin
        s1_req_addr <= T_2319;
      end
    end
    if(1'h0) begin
    end else begin
      if(metaReadArb_io_out_valid) begin
        s1_req_tag <= io_cpu_req_bits_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(metaReadArb_io_out_valid) begin
        s1_req_cmd <= io_cpu_req_bits_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(metaReadArb_io_out_valid) begin
        s1_req_typ <= io_cpu_req_bits_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(metaReadArb_io_out_valid) begin
        s1_req_phys <= io_cpu_req_bits_phys;
      end
    end
    if(1'h0) begin
    end else begin
      if(metaReadArb_io_out_valid) begin
        s1_req_data <= io_cpu_req_bits_data;
      end
    end
    if(1'h0) begin
    end else begin
      s1_flush_valid <= T_4530;
    end
    if(reset) begin
      grant_wait <= 1'h0;
    end else begin
      if(T_3776) begin
        grant_wait <= 1'h0;
      end else begin
        if(T_3741) begin
          grant_wait <= 1'h1;
        end
      end
    end
    if(reset) begin
      release_ack_wait <= 1'h0;
    end else begin
      if(T_4410) begin
        if(releaseDone) begin
          release_ack_wait <= 1'h1;
        end else begin
          if(io_mem_grant_valid) begin
            if(grantIsVoluntary) begin
              release_ack_wait <= 1'h0;
            end
          end
        end
      end else begin
        if(io_mem_grant_valid) begin
          if(grantIsVoluntary) begin
            release_ack_wait <= 1'h0;
          end
        end
      end
    end
    if(reset) begin
      release_state <= 3'h0;
    end else begin
      if(T_4437) begin
        release_state <= 3'h0;
      end else begin
        if(T_4410) begin
          if(releaseDone) begin
            release_state <= 3'h6;
          end else begin
            if(T_4407) begin
              if(releaseDone) begin
                release_state <= 3'h7;
              end else begin
                if(releaseDone) begin
                  release_state <= 3'h0;
                end else begin
                  if(s2_probe) begin
                    if(T_4399) begin
                      release_state <= 3'h5;
                    end else begin
                      if(T_4394) begin
                        release_state <= 3'h4;
                      end else begin
                        if(T_4221) begin
                          release_state <= 3'h3;
                        end else begin
                          if(T_4381) begin
                            release_state <= 3'h2;
                          end
                        end
                      end
                    end
                  end else begin
                    if(T_4381) begin
                      release_state <= 3'h2;
                    end
                  end
                end
              end
            end else begin
              if(releaseDone) begin
                release_state <= 3'h0;
              end else begin
                if(s2_probe) begin
                  if(T_4399) begin
                    release_state <= 3'h5;
                  end else begin
                    if(T_4394) begin
                      release_state <= 3'h4;
                    end else begin
                      if(T_4221) begin
                        release_state <= 3'h3;
                      end else begin
                        if(T_4381) begin
                          release_state <= 3'h2;
                        end
                      end
                    end
                  end
                end else begin
                  if(T_4381) begin
                    release_state <= 3'h2;
                  end
                end
              end
            end
          end
        end else begin
          if(T_4407) begin
            if(releaseDone) begin
              release_state <= 3'h7;
            end else begin
              if(releaseDone) begin
                release_state <= 3'h0;
              end else begin
                if(s2_probe) begin
                  if(T_4399) begin
                    release_state <= 3'h5;
                  end else begin
                    if(T_4394) begin
                      release_state <= 3'h4;
                    end else begin
                      if(T_4221) begin
                        release_state <= 3'h3;
                      end else begin
                        release_state <= GEN_77;
                      end
                    end
                  end
                end else begin
                  release_state <= GEN_77;
                end
              end
            end
          end else begin
            if(releaseDone) begin
              release_state <= 3'h0;
            end else begin
              if(s2_probe) begin
                if(T_4399) begin
                  release_state <= 3'h5;
                end else begin
                  if(T_4394) begin
                    release_state <= 3'h4;
                  end else begin
                    if(T_4221) begin
                      release_state <= 3'h3;
                    end else begin
                      release_state <= GEN_77;
                    end
                  end
                end
              end else begin
                release_state <= GEN_77;
              end
            end
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      pstore2_valid <= T_3011;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= s1_valid_masked;
    end
    if(reset) begin
      s2_probe <= 1'h0;
    end else begin
      s2_probe <= s1_probe;
    end
    if(1'h0) begin
    end else begin
      T_2500 <= T_2249;
    end
    if(1'h0) begin
    end else begin
      if(T_2568) begin
        s2_req_addr <= s1_paddr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2568) begin
        s2_req_tag <= s1_req_tag;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2568) begin
        s2_req_cmd <= s1_req_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2568) begin
        s2_req_typ <= s1_req_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2568) begin
        s2_req_phys <= s1_req_phys;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2568) begin
        s2_req_data <= s1_req_data;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2568) begin
        s2_uncached <= T_2570;
      end
    end
    if(1'h0) begin
    end else begin
      s2_flush_valid <= s1_flush_valid;
    end
    if(1'h0) begin
    end else begin
      if(io_mem_grant_valid) begin
        if(grantIsUncached) begin
          s2_data <= io_mem_grant_bits_data;
        end else begin
          if(T_2585) begin
            s2_data <= data_io_resp_0;
          end
        end
      end else begin
        if(T_2585) begin
          s2_data <= data_io_resp_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_probe) begin
        s2_probe_way <= s1_hit_way;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_probe) begin
        s2_probe_state_state <= s1_hit_state_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_valid_not_nacked) begin
        s2_hit_way <= s1_hit_way;
      end
    end
    if(1'h0) begin
    end else begin
      if(s1_valid_not_nacked) begin
        s2_hit_state_state <= s1_hit_state_state;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2568) begin
        T_2663 <= s1_victim_way;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2568) begin
        s2_victim_tag <= GEN_0;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2568) begin
        T_2839_state <= GEN_1;
      end
    end
    if(1'h0) begin
    end else begin
      T_2910 <= T_2909;
    end
    if(reset) begin
      lrscCount <= 5'h0;
    end else begin
      if(io_cpu_invalidate_lr) begin
        lrscCount <= 5'h0;
      end else begin
        if(lrscValid) begin
          lrscCount <= T_2934;
        end
      end
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      if(T_2938) begin
        pstore1_cmd <= s1_req_cmd;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2938) begin
        pstore1_typ <= s1_req_typ;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2938) begin
        pstore1_addr <= s1_paddr;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2938) begin
        pstore1_data <= io_cpu_s1_data;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2938) begin
        pstore1_way <= s1_hit_way;
      end
    end
    if(1'h0) begin
    end else begin
      T_2992 <= T_3005;
    end
    if(1'h0) begin
    end else begin
      if(advance_pstore1) begin
        pstore2_addr <= pstore1_addr;
      end
    end
    if(1'h0) begin
    end else begin
      if(advance_pstore1) begin
        pstore2_way <= pstore1_way;
      end
    end
    if(1'h0) begin
    end else begin
      if(advance_pstore1) begin
        pstore2_storegen_data <= pstore1_storegen_data;
      end
    end
    if(1'h0) begin
    end else begin
      if(advance_pstore1) begin
        pstore2_storegen_mask <= T_3038;
      end
    end
    if(reset) begin
      refillCount <= 3'h0;
    end else begin
      if(T_3768) begin
        refillCount <= T_3774;
      end
    end
    if(reset) begin
      writebackCount <= 3'h0;
    end else begin
      if(T_3936) begin
        writebackCount <= T_3942;
      end
    end
    if(1'h0) begin
    end else begin
      s1_release_data_valid <= T_3949;
    end
    if(1'h0) begin
    end else begin
      s2_release_data_valid <= T_3952;
    end
    if(1'h0) begin
    end else begin
      doUncachedResp <= io_cpu_replay_next;
    end
    if(reset) begin
      flushed <= 1'h1;
    end else begin
      if(flushing) begin
        if(s2_flush_valid) begin
          if(T_4535) begin
            flushed <= 1'h1;
          end else begin
            if(T_3741) begin
              flushed <= 1'h0;
            end
          end
        end else begin
          if(T_3741) begin
            flushed <= 1'h0;
          end
        end
      end else begin
        if(T_3741) begin
          flushed <= 1'h0;
        end
      end
    end
    if(reset) begin
      flushing <= 1'h0;
    end else begin
      if(flushing) begin
        if(T_4544) begin
          flushing <= 1'h0;
        end else begin
          if(T_4512) begin
            if(T_4514) begin
              flushing <= T_2655;
            end
          end
        end
      end else begin
        if(T_4512) begin
          if(T_4514) begin
            flushing <= T_2655;
          end
        end
      end
    end
    if(reset) begin
      T_4508 <= 7'h0;
    end else begin
      if(flushing) begin
        if(s2_flush_valid) begin
          T_4508 <= T_4538;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_2916) begin
          $fwrite(32'h80000002,"Assertion failed: DCache exception occurred - cache response not killed.\n    at dcache.scala:167 assert(!(Reg(next=\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_2916) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_3000) begin
          $fwrite(32'h80000002,"Assertion failed\n    at dcache.scala:204 assert(!s2_store_valid || !pstore1_held)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_3000) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (s2_uncached & T_3740) begin
          $fwrite(32'h80000002,"Assertion failed: cache hit on uncached access\n    at dcache.scala:267 assert(!s2_valid_masked || !s2_hit_state.isValid(), ---cache hit on uncached access---)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (s2_uncached & T_3740) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_mem_grant_valid & T_3765) begin
          $fwrite(32'h80000002,"Assertion failed: unexpected grant\n    at dcache.scala:283 assert(grant_wait || grantIsVoluntary && release_ack_wait, ---unexpected grant---)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_mem_grant_valid & T_3765) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_3785) begin
          $fwrite(32'h80000002,"Assertion failed\n    at dcache.scala:294 assert(dataArb.io.in(1).ready || !dataArb.io.in(1).valid)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_3785) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_3797) begin
          $fwrite(32'h80000002,"Assertion failed\n    at dcache.scala:302 assert(!metaWriteArb.io.in(1).valid || metaWriteArb.io.in(1).ready)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_3797) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (fq_io_enq_valid & T_3916) begin
          $fwrite(32'h80000002,"Assertion failed\n    at dcache.scala:312 when (fq.io.enq.valid) { assert(fq.io.enq.ready) }\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (fq_io_enq_valid & T_3916) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_4381 & T_4387) begin
          $fwrite(32'h80000002,"Assertion failed\n    at dcache.scala:338 assert(!s2_hit_state.isValid())\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_4381 & T_4387) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (doUncachedResp & T_4448) begin
          $fwrite(32'h80000002,"Assertion failed\n    at dcache.scala:395 assert(!s2_valid_hit)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (doUncachedResp & T_4448) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_4504) begin
          $fwrite(32'h80000002,"Assertion failed: unsupported D$ operation\n    at dcache.scala:418 assert(!(s1_valid_masked && s1_read && s1_write), ---unsupported D$ operation---)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_4504) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module ClientUncachedTileLinkIOArbiter(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input   io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output  io_in_0_grant_bits_client_xact_id,
  output [1:0] io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_acquire_ready,
  output  io_out_acquire_valid,
  output [25:0] io_out_acquire_bits_addr_block,
  output  io_out_acquire_bits_client_xact_id,
  output [2:0] io_out_acquire_bits_addr_beat,
  output  io_out_acquire_bits_is_builtin_type,
  output [2:0] io_out_acquire_bits_a_type,
  output [11:0] io_out_acquire_bits_union,
  output [63:0] io_out_acquire_bits_data,
  output  io_out_grant_ready,
  input   io_out_grant_valid,
  input  [2:0] io_out_grant_bits_addr_beat,
  input   io_out_grant_bits_client_xact_id,
  input  [1:0] io_out_grant_bits_manager_xact_id,
  input   io_out_grant_bits_is_builtin_type,
  input  [3:0] io_out_grant_bits_g_type,
  input  [63:0] io_out_grant_bits_data
);
  assign io_in_0_acquire_ready = io_out_acquire_ready;
  assign io_in_0_grant_valid = io_out_grant_valid;
  assign io_in_0_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_0_grant_bits_data = io_out_grant_bits_data;
  assign io_out_acquire_valid = io_in_0_acquire_valid;
  assign io_out_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign io_out_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign io_out_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign io_out_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign io_out_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign io_out_acquire_bits_union = io_in_0_acquire_bits_union;
  assign io_out_acquire_bits_data = io_in_0_acquire_bits_data;
  assign io_out_grant_ready = io_in_0_grant_ready;
endmodule
module HellaCacheArbiter(
  input   clk,
  input   reset,
  output  io_requestor_0_req_ready,
  input   io_requestor_0_req_valid,
  input  [31:0] io_requestor_0_req_bits_addr,
  input  [8:0] io_requestor_0_req_bits_tag,
  input  [4:0] io_requestor_0_req_bits_cmd,
  input  [2:0] io_requestor_0_req_bits_typ,
  input   io_requestor_0_req_bits_phys,
  input  [31:0] io_requestor_0_req_bits_data,
  input   io_requestor_0_s1_kill,
  input  [31:0] io_requestor_0_s1_data,
  output  io_requestor_0_s2_nack,
  output  io_requestor_0_resp_valid,
  output [31:0] io_requestor_0_resp_bits_addr,
  output [8:0] io_requestor_0_resp_bits_tag,
  output [4:0] io_requestor_0_resp_bits_cmd,
  output [2:0] io_requestor_0_resp_bits_typ,
  output [31:0] io_requestor_0_resp_bits_data,
  output  io_requestor_0_resp_bits_replay,
  output  io_requestor_0_resp_bits_has_data,
  output [31:0] io_requestor_0_resp_bits_data_word_bypass,
  output [31:0] io_requestor_0_resp_bits_store_data,
  output  io_requestor_0_replay_next,
  output  io_requestor_0_xcpt_ma_ld,
  output  io_requestor_0_xcpt_ma_st,
  output  io_requestor_0_xcpt_pf_ld,
  output  io_requestor_0_xcpt_pf_st,
  input   io_requestor_0_invalidate_lr,
  output  io_requestor_0_ordered,
  input   io_mem_req_ready,
  output  io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [8:0] io_mem_req_bits_tag,
  output [4:0] io_mem_req_bits_cmd,
  output [2:0] io_mem_req_bits_typ,
  output  io_mem_req_bits_phys,
  output [31:0] io_mem_req_bits_data,
  output  io_mem_s1_kill,
  output [31:0] io_mem_s1_data,
  input   io_mem_s2_nack,
  input   io_mem_resp_valid,
  input  [31:0] io_mem_resp_bits_addr,
  input  [8:0] io_mem_resp_bits_tag,
  input  [4:0] io_mem_resp_bits_cmd,
  input  [2:0] io_mem_resp_bits_typ,
  input  [31:0] io_mem_resp_bits_data,
  input   io_mem_resp_bits_replay,
  input   io_mem_resp_bits_has_data,
  input  [31:0] io_mem_resp_bits_data_word_bypass,
  input  [31:0] io_mem_resp_bits_store_data,
  input   io_mem_replay_next,
  input   io_mem_xcpt_ma_ld,
  input   io_mem_xcpt_ma_st,
  input   io_mem_xcpt_pf_ld,
  input   io_mem_xcpt_pf_st,
  output  io_mem_invalidate_lr,
  input   io_mem_ordered
);
  assign io_requestor_0_req_ready = io_mem_req_ready;
  assign io_requestor_0_s2_nack = io_mem_s2_nack;
  assign io_requestor_0_resp_valid = io_mem_resp_valid;
  assign io_requestor_0_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_0_resp_bits_tag = io_mem_resp_bits_tag;
  assign io_requestor_0_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_0_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_0_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_0_resp_bits_replay = io_mem_resp_bits_replay;
  assign io_requestor_0_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_0_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass;
  assign io_requestor_0_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_0_replay_next = io_mem_replay_next;
  assign io_requestor_0_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_0_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_0_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_0_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_0_ordered = io_mem_ordered;
  assign io_mem_req_valid = io_requestor_0_req_valid;
  assign io_mem_req_bits_addr = io_requestor_0_req_bits_addr;
  assign io_mem_req_bits_tag = io_requestor_0_req_bits_tag;
  assign io_mem_req_bits_cmd = io_requestor_0_req_bits_cmd;
  assign io_mem_req_bits_typ = io_requestor_0_req_bits_typ;
  assign io_mem_req_bits_phys = io_requestor_0_req_bits_phys;
  assign io_mem_req_bits_data = io_requestor_0_req_bits_data;
  assign io_mem_s1_kill = io_requestor_0_s1_kill;
  assign io_mem_s1_data = io_requestor_0_s1_data;
  assign io_mem_invalidate_lr = io_requestor_0_invalidate_lr;
endmodule
module RocketTile(
  input   clk,
  input   reset,
  input   io_cached_0_acquire_ready,
  output  io_cached_0_acquire_valid,
  output [25:0] io_cached_0_acquire_bits_addr_block,
  output  io_cached_0_acquire_bits_client_xact_id,
  output [2:0] io_cached_0_acquire_bits_addr_beat,
  output  io_cached_0_acquire_bits_is_builtin_type,
  output [2:0] io_cached_0_acquire_bits_a_type,
  output [11:0] io_cached_0_acquire_bits_union,
  output [63:0] io_cached_0_acquire_bits_data,
  output  io_cached_0_probe_ready,
  input   io_cached_0_probe_valid,
  input  [25:0] io_cached_0_probe_bits_addr_block,
  input  [1:0] io_cached_0_probe_bits_p_type,
  input   io_cached_0_release_ready,
  output  io_cached_0_release_valid,
  output [2:0] io_cached_0_release_bits_addr_beat,
  output [25:0] io_cached_0_release_bits_addr_block,
  output  io_cached_0_release_bits_client_xact_id,
  output  io_cached_0_release_bits_voluntary,
  output [2:0] io_cached_0_release_bits_r_type,
  output [63:0] io_cached_0_release_bits_data,
  output  io_cached_0_grant_ready,
  input   io_cached_0_grant_valid,
  input  [2:0] io_cached_0_grant_bits_addr_beat,
  input   io_cached_0_grant_bits_client_xact_id,
  input  [1:0] io_cached_0_grant_bits_manager_xact_id,
  input   io_cached_0_grant_bits_is_builtin_type,
  input  [3:0] io_cached_0_grant_bits_g_type,
  input  [63:0] io_cached_0_grant_bits_data,
  input   io_cached_0_grant_bits_manager_id,
  input   io_cached_0_finish_ready,
  output  io_cached_0_finish_valid,
  output [1:0] io_cached_0_finish_bits_manager_xact_id,
  output  io_cached_0_finish_bits_manager_id,
  input   io_uncached_0_acquire_ready,
  output  io_uncached_0_acquire_valid,
  output [25:0] io_uncached_0_acquire_bits_addr_block,
  output  io_uncached_0_acquire_bits_client_xact_id,
  output [2:0] io_uncached_0_acquire_bits_addr_beat,
  output  io_uncached_0_acquire_bits_is_builtin_type,
  output [2:0] io_uncached_0_acquire_bits_a_type,
  output [11:0] io_uncached_0_acquire_bits_union,
  output [63:0] io_uncached_0_acquire_bits_data,
  output  io_uncached_0_grant_ready,
  input   io_uncached_0_grant_valid,
  input  [2:0] io_uncached_0_grant_bits_addr_beat,
  input   io_uncached_0_grant_bits_client_xact_id,
  input  [1:0] io_uncached_0_grant_bits_manager_xact_id,
  input   io_uncached_0_grant_bits_is_builtin_type,
  input  [3:0] io_uncached_0_grant_bits_g_type,
  input  [63:0] io_uncached_0_grant_bits_data,
  input   io_prci_reset,
  input   io_prci_id,
  input   io_prci_interrupts_meip,
  input   io_prci_interrupts_seip,
  input   io_prci_interrupts_debug,
  input   io_prci_interrupts_mtip,
  input   io_prci_interrupts_msip
);
//<CJ> RESET_VECTOR_ADDR
  parameter RESET_VECTOR_ADDR = 60000000;

  wire  core_clk;
  wire  core_reset;
  wire  core_io_prci_reset;
  wire  core_io_prci_id;
  wire  core_io_prci_interrupts_meip;
  wire  core_io_prci_interrupts_seip;
  wire  core_io_prci_interrupts_debug;
  wire  core_io_prci_interrupts_mtip;
  wire  core_io_prci_interrupts_msip;
  wire  core_io_imem_req_valid;
  wire [31:0] core_io_imem_req_bits_pc;
  wire  core_io_imem_req_bits_speculative;
  wire  core_io_imem_resp_ready;
  wire  core_io_imem_resp_valid;
  wire [31:0] core_io_imem_resp_bits_pc;
  wire [31:0] core_io_imem_resp_bits_data_0;
  wire  core_io_imem_resp_bits_mask;
  wire  core_io_imem_resp_bits_xcpt_if;
  wire  core_io_imem_resp_bits_replay;
  wire  core_io_imem_btb_resp_valid;
  wire  core_io_imem_btb_resp_bits_taken;
  wire  core_io_imem_btb_resp_bits_mask;
  wire  core_io_imem_btb_resp_bits_bridx;
  wire [31:0] core_io_imem_btb_resp_bits_target;
  wire  core_io_imem_btb_resp_bits_entry;
  wire  core_io_imem_btb_resp_bits_bht_history;
  wire [1:0] core_io_imem_btb_resp_bits_bht_value;
  wire  core_io_imem_btb_update_valid;
  wire  core_io_imem_btb_update_bits_prediction_valid;
  wire  core_io_imem_btb_update_bits_prediction_bits_taken;
  wire  core_io_imem_btb_update_bits_prediction_bits_mask;
  wire  core_io_imem_btb_update_bits_prediction_bits_bridx;
  wire [31:0] core_io_imem_btb_update_bits_prediction_bits_target;
  wire  core_io_imem_btb_update_bits_prediction_bits_entry;
  wire  core_io_imem_btb_update_bits_prediction_bits_bht_history;
  wire [1:0] core_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire [31:0] core_io_imem_btb_update_bits_pc;
  wire [31:0] core_io_imem_btb_update_bits_target;
  wire  core_io_imem_btb_update_bits_taken;
  wire  core_io_imem_btb_update_bits_isJump;
  wire  core_io_imem_btb_update_bits_isReturn;
  wire [31:0] core_io_imem_btb_update_bits_br_pc;
  wire  core_io_imem_bht_update_valid;
  wire  core_io_imem_bht_update_bits_prediction_valid;
  wire  core_io_imem_bht_update_bits_prediction_bits_taken;
  wire  core_io_imem_bht_update_bits_prediction_bits_mask;
  wire  core_io_imem_bht_update_bits_prediction_bits_bridx;
  wire [31:0] core_io_imem_bht_update_bits_prediction_bits_target;
  wire  core_io_imem_bht_update_bits_prediction_bits_entry;
  wire  core_io_imem_bht_update_bits_prediction_bits_bht_history;
  wire [1:0] core_io_imem_bht_update_bits_prediction_bits_bht_value;
  wire [31:0] core_io_imem_bht_update_bits_pc;
  wire  core_io_imem_bht_update_bits_taken;
  wire  core_io_imem_bht_update_bits_mispredict;
  wire  core_io_imem_ras_update_valid;
  wire  core_io_imem_ras_update_bits_isCall;
  wire  core_io_imem_ras_update_bits_isReturn;
  wire [31:0] core_io_imem_ras_update_bits_returnAddr;
  wire  core_io_imem_ras_update_bits_prediction_valid;
  wire  core_io_imem_ras_update_bits_prediction_bits_taken;
  wire  core_io_imem_ras_update_bits_prediction_bits_mask;
  wire  core_io_imem_ras_update_bits_prediction_bits_bridx;
  wire [31:0] core_io_imem_ras_update_bits_prediction_bits_target;
  wire  core_io_imem_ras_update_bits_prediction_bits_entry;
  wire  core_io_imem_ras_update_bits_prediction_bits_bht_history;
  wire [1:0] core_io_imem_ras_update_bits_prediction_bits_bht_value;
  wire  core_io_imem_flush_icache;
  wire  core_io_imem_flush_tlb;
  wire [31:0] core_io_imem_npc;
  wire  core_io_dmem_req_ready;
  wire  core_io_dmem_req_valid;
  wire [31:0] core_io_dmem_req_bits_addr;
  wire [8:0] core_io_dmem_req_bits_tag;
  wire [4:0] core_io_dmem_req_bits_cmd;
  wire [2:0] core_io_dmem_req_bits_typ;
  wire  core_io_dmem_req_bits_phys;
  wire [31:0] core_io_dmem_req_bits_data;
  wire  core_io_dmem_s1_kill;
  wire [31:0] core_io_dmem_s1_data;
  wire  core_io_dmem_s2_nack;
  wire  core_io_dmem_resp_valid;
  wire [31:0] core_io_dmem_resp_bits_addr;
  wire [8:0] core_io_dmem_resp_bits_tag;
  wire [4:0] core_io_dmem_resp_bits_cmd;
  wire [2:0] core_io_dmem_resp_bits_typ;
  wire [31:0] core_io_dmem_resp_bits_data;
  wire  core_io_dmem_resp_bits_replay;
  wire  core_io_dmem_resp_bits_has_data;
  wire [31:0] core_io_dmem_resp_bits_data_word_bypass;
  wire [31:0] core_io_dmem_resp_bits_store_data;
  wire  core_io_dmem_replay_next;
  wire  core_io_dmem_xcpt_ma_ld;
  wire  core_io_dmem_xcpt_ma_st;
  wire  core_io_dmem_xcpt_pf_ld;
  wire  core_io_dmem_xcpt_pf_st;
  wire  core_io_dmem_invalidate_lr;
  wire  core_io_dmem_ordered;
  wire [6:0] core_io_ptw_ptbr_asid;
  wire [21:0] core_io_ptw_ptbr_ppn;
  wire  core_io_ptw_invalidate;
  wire  core_io_ptw_status_debug;
  wire [1:0] core_io_ptw_status_prv;
  wire  core_io_ptw_status_sd;
  wire [30:0] core_io_ptw_status_zero3;
  wire  core_io_ptw_status_sd_rv32;
  wire [1:0] core_io_ptw_status_zero2;
  wire [4:0] core_io_ptw_status_vm;
  wire [3:0] core_io_ptw_status_zero1;
  wire  core_io_ptw_status_mxr;
  wire  core_io_ptw_status_pum;
  wire  core_io_ptw_status_mprv;
  wire [1:0] core_io_ptw_status_xs;
  wire [1:0] core_io_ptw_status_fs;
  wire [1:0] core_io_ptw_status_mpp;
  wire [1:0] core_io_ptw_status_hpp;
  wire  core_io_ptw_status_spp;
  wire  core_io_ptw_status_mpie;
  wire  core_io_ptw_status_hpie;
  wire  core_io_ptw_status_spie;
  wire  core_io_ptw_status_upie;
  wire  core_io_ptw_status_mie;
  wire  core_io_ptw_status_hie;
  wire  core_io_ptw_status_sie;
  wire  core_io_ptw_status_uie;
  wire [31:0] core_io_fpu_inst;
  wire [31:0] core_io_fpu_fromint_data;
  wire [2:0] core_io_fpu_fcsr_rm;
  wire  core_io_fpu_fcsr_flags_valid;
  wire [4:0] core_io_fpu_fcsr_flags_bits;
  wire [63:0] core_io_fpu_store_data;
  wire [31:0] core_io_fpu_toint_data;
  wire  core_io_fpu_dmem_resp_val;
  wire [2:0] core_io_fpu_dmem_resp_type;
  wire [4:0] core_io_fpu_dmem_resp_tag;
  wire [63:0] core_io_fpu_dmem_resp_data;
  wire  core_io_fpu_valid;
  wire  core_io_fpu_fcsr_rdy;
  wire  core_io_fpu_nack_mem;
  wire  core_io_fpu_illegal_rm;
  wire  core_io_fpu_killx;
  wire  core_io_fpu_killm;
  wire [4:0] core_io_fpu_dec_cmd;
  wire  core_io_fpu_dec_ldst;
  wire  core_io_fpu_dec_wen;
  wire  core_io_fpu_dec_ren1;
  wire  core_io_fpu_dec_ren2;
  wire  core_io_fpu_dec_ren3;
  wire  core_io_fpu_dec_swap12;
  wire  core_io_fpu_dec_swap23;
  wire  core_io_fpu_dec_single;
  wire  core_io_fpu_dec_fromint;
  wire  core_io_fpu_dec_toint;
  wire  core_io_fpu_dec_fastpipe;
  wire  core_io_fpu_dec_fma;
  wire  core_io_fpu_dec_div;
  wire  core_io_fpu_dec_sqrt;
  wire  core_io_fpu_dec_round;
  wire  core_io_fpu_dec_wflags;
  wire  core_io_fpu_sboard_set;
  wire  core_io_fpu_sboard_clr;
  wire [4:0] core_io_fpu_sboard_clra;
  wire  core_io_fpu_cp_req_ready;
  wire  core_io_fpu_cp_req_valid;
  wire [4:0] core_io_fpu_cp_req_bits_cmd;
  wire  core_io_fpu_cp_req_bits_ldst;
  wire  core_io_fpu_cp_req_bits_wen;
  wire  core_io_fpu_cp_req_bits_ren1;
  wire  core_io_fpu_cp_req_bits_ren2;
  wire  core_io_fpu_cp_req_bits_ren3;
  wire  core_io_fpu_cp_req_bits_swap12;
  wire  core_io_fpu_cp_req_bits_swap23;
  wire  core_io_fpu_cp_req_bits_single;
  wire  core_io_fpu_cp_req_bits_fromint;
  wire  core_io_fpu_cp_req_bits_toint;
  wire  core_io_fpu_cp_req_bits_fastpipe;
  wire  core_io_fpu_cp_req_bits_fma;
  wire  core_io_fpu_cp_req_bits_div;
  wire  core_io_fpu_cp_req_bits_sqrt;
  wire  core_io_fpu_cp_req_bits_round;
  wire  core_io_fpu_cp_req_bits_wflags;
  wire [2:0] core_io_fpu_cp_req_bits_rm;
  wire [1:0] core_io_fpu_cp_req_bits_typ;
  wire [64:0] core_io_fpu_cp_req_bits_in1;
  wire [64:0] core_io_fpu_cp_req_bits_in2;
  wire [64:0] core_io_fpu_cp_req_bits_in3;
  wire  core_io_fpu_cp_resp_ready;
  wire  core_io_fpu_cp_resp_valid;
  wire [64:0] core_io_fpu_cp_resp_bits_data;
  wire [4:0] core_io_fpu_cp_resp_bits_exc;
  wire  core_io_rocc_cmd_ready;
  wire  core_io_rocc_cmd_valid;
  wire [6:0] core_io_rocc_cmd_bits_inst_funct;
  wire [4:0] core_io_rocc_cmd_bits_inst_rs2;
  wire [4:0] core_io_rocc_cmd_bits_inst_rs1;
  wire  core_io_rocc_cmd_bits_inst_xd;
  wire  core_io_rocc_cmd_bits_inst_xs1;
  wire  core_io_rocc_cmd_bits_inst_xs2;
  wire [4:0] core_io_rocc_cmd_bits_inst_rd;
  wire [6:0] core_io_rocc_cmd_bits_inst_opcode;
  wire [31:0] core_io_rocc_cmd_bits_rs1;
  wire [31:0] core_io_rocc_cmd_bits_rs2;
  wire  core_io_rocc_cmd_bits_status_debug;
  wire [1:0] core_io_rocc_cmd_bits_status_prv;
  wire  core_io_rocc_cmd_bits_status_sd;
  wire [30:0] core_io_rocc_cmd_bits_status_zero3;
  wire  core_io_rocc_cmd_bits_status_sd_rv32;
  wire [1:0] core_io_rocc_cmd_bits_status_zero2;
  wire [4:0] core_io_rocc_cmd_bits_status_vm;
  wire [3:0] core_io_rocc_cmd_bits_status_zero1;
  wire  core_io_rocc_cmd_bits_status_mxr;
  wire  core_io_rocc_cmd_bits_status_pum;
  wire  core_io_rocc_cmd_bits_status_mprv;
  wire [1:0] core_io_rocc_cmd_bits_status_xs;
  wire [1:0] core_io_rocc_cmd_bits_status_fs;
  wire [1:0] core_io_rocc_cmd_bits_status_mpp;
  wire [1:0] core_io_rocc_cmd_bits_status_hpp;
  wire  core_io_rocc_cmd_bits_status_spp;
  wire  core_io_rocc_cmd_bits_status_mpie;
  wire  core_io_rocc_cmd_bits_status_hpie;
  wire  core_io_rocc_cmd_bits_status_spie;
  wire  core_io_rocc_cmd_bits_status_upie;
  wire  core_io_rocc_cmd_bits_status_mie;
  wire  core_io_rocc_cmd_bits_status_hie;
  wire  core_io_rocc_cmd_bits_status_sie;
  wire  core_io_rocc_cmd_bits_status_uie;
  wire  core_io_rocc_resp_ready;
  wire  core_io_rocc_resp_valid;
  wire [4:0] core_io_rocc_resp_bits_rd;
  wire [31:0] core_io_rocc_resp_bits_data;
  wire  core_io_rocc_mem_req_ready;
  wire  core_io_rocc_mem_req_valid;
  wire [31:0] core_io_rocc_mem_req_bits_addr;
  wire [8:0] core_io_rocc_mem_req_bits_tag;
  wire [4:0] core_io_rocc_mem_req_bits_cmd;
  wire [2:0] core_io_rocc_mem_req_bits_typ;
  wire  core_io_rocc_mem_req_bits_phys;
  wire [31:0] core_io_rocc_mem_req_bits_data;
  wire  core_io_rocc_mem_s1_kill;
  wire [31:0] core_io_rocc_mem_s1_data;
  wire  core_io_rocc_mem_s2_nack;
  wire  core_io_rocc_mem_resp_valid;
  wire [31:0] core_io_rocc_mem_resp_bits_addr;
  wire [8:0] core_io_rocc_mem_resp_bits_tag;
  wire [4:0] core_io_rocc_mem_resp_bits_cmd;
  wire [2:0] core_io_rocc_mem_resp_bits_typ;
  wire [31:0] core_io_rocc_mem_resp_bits_data;
  wire  core_io_rocc_mem_resp_bits_replay;
  wire  core_io_rocc_mem_resp_bits_has_data;
  wire [31:0] core_io_rocc_mem_resp_bits_data_word_bypass;
  wire [31:0] core_io_rocc_mem_resp_bits_store_data;
  wire  core_io_rocc_mem_replay_next;
  wire  core_io_rocc_mem_xcpt_ma_ld;
  wire  core_io_rocc_mem_xcpt_ma_st;
  wire  core_io_rocc_mem_xcpt_pf_ld;
  wire  core_io_rocc_mem_xcpt_pf_st;
  wire  core_io_rocc_mem_invalidate_lr;
  wire  core_io_rocc_mem_ordered;
  wire  core_io_rocc_busy;
  wire  core_io_rocc_interrupt;
  wire  core_io_rocc_autl_acquire_ready;
  wire  core_io_rocc_autl_acquire_valid;
  wire [25:0] core_io_rocc_autl_acquire_bits_addr_block;
  wire  core_io_rocc_autl_acquire_bits_client_xact_id;
  wire [2:0] core_io_rocc_autl_acquire_bits_addr_beat;
  wire  core_io_rocc_autl_acquire_bits_is_builtin_type;
  wire [2:0] core_io_rocc_autl_acquire_bits_a_type;
  wire [11:0] core_io_rocc_autl_acquire_bits_union;
  wire [63:0] core_io_rocc_autl_acquire_bits_data;
  wire  core_io_rocc_autl_grant_ready;
  wire  core_io_rocc_autl_grant_valid;
  wire [2:0] core_io_rocc_autl_grant_bits_addr_beat;
  wire  core_io_rocc_autl_grant_bits_client_xact_id;
  wire [1:0] core_io_rocc_autl_grant_bits_manager_xact_id;
  wire  core_io_rocc_autl_grant_bits_is_builtin_type;
  wire [3:0] core_io_rocc_autl_grant_bits_g_type;
  wire [63:0] core_io_rocc_autl_grant_bits_data;
  wire  core_io_rocc_fpu_req_ready;
  wire  core_io_rocc_fpu_req_valid;
  wire [4:0] core_io_rocc_fpu_req_bits_cmd;
  wire  core_io_rocc_fpu_req_bits_ldst;
  wire  core_io_rocc_fpu_req_bits_wen;
  wire  core_io_rocc_fpu_req_bits_ren1;
  wire  core_io_rocc_fpu_req_bits_ren2;
  wire  core_io_rocc_fpu_req_bits_ren3;
  wire  core_io_rocc_fpu_req_bits_swap12;
  wire  core_io_rocc_fpu_req_bits_swap23;
  wire  core_io_rocc_fpu_req_bits_single;
  wire  core_io_rocc_fpu_req_bits_fromint;
  wire  core_io_rocc_fpu_req_bits_toint;
  wire  core_io_rocc_fpu_req_bits_fastpipe;
  wire  core_io_rocc_fpu_req_bits_fma;
  wire  core_io_rocc_fpu_req_bits_div;
  wire  core_io_rocc_fpu_req_bits_sqrt;
  wire  core_io_rocc_fpu_req_bits_round;
  wire  core_io_rocc_fpu_req_bits_wflags;
  wire [2:0] core_io_rocc_fpu_req_bits_rm;
  wire [1:0] core_io_rocc_fpu_req_bits_typ;
  wire [64:0] core_io_rocc_fpu_req_bits_in1;
  wire [64:0] core_io_rocc_fpu_req_bits_in2;
  wire [64:0] core_io_rocc_fpu_req_bits_in3;
  wire  core_io_rocc_fpu_resp_ready;
  wire  core_io_rocc_fpu_resp_valid;
  wire [64:0] core_io_rocc_fpu_resp_bits_data;
  wire [4:0] core_io_rocc_fpu_resp_bits_exc;
  wire  core_io_rocc_exception;
  wire [11:0] core_io_rocc_csr_waddr;
  wire [31:0] core_io_rocc_csr_wdata;
  wire  core_io_rocc_csr_wen;
  wire  core_io_rocc_host_id;
  wire  icache_clk;
  wire  icache_reset;
  wire  icache_io_cpu_req_valid;
  wire [31:0] icache_io_cpu_req_bits_pc;
  wire  icache_io_cpu_req_bits_speculative;
  wire  icache_io_cpu_resp_ready;
  wire  icache_io_cpu_resp_valid;
  wire [31:0] icache_io_cpu_resp_bits_pc;
  wire [31:0] icache_io_cpu_resp_bits_data_0;
  wire  icache_io_cpu_resp_bits_mask;
  wire  icache_io_cpu_resp_bits_xcpt_if;
  wire  icache_io_cpu_resp_bits_replay;
  wire  icache_io_cpu_btb_resp_valid;
  wire  icache_io_cpu_btb_resp_bits_taken;
  wire  icache_io_cpu_btb_resp_bits_mask;
  wire  icache_io_cpu_btb_resp_bits_bridx;
  wire [31:0] icache_io_cpu_btb_resp_bits_target;
  wire  icache_io_cpu_btb_resp_bits_entry;
  wire  icache_io_cpu_btb_resp_bits_bht_history;
  wire [1:0] icache_io_cpu_btb_resp_bits_bht_value;
  wire  icache_io_cpu_btb_update_valid;
  wire  icache_io_cpu_btb_update_bits_prediction_valid;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_taken;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_mask;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_bridx;
  wire [31:0] icache_io_cpu_btb_update_bits_prediction_bits_target;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_entry;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_bht_history;
  wire [1:0] icache_io_cpu_btb_update_bits_prediction_bits_bht_value;
  wire [31:0] icache_io_cpu_btb_update_bits_pc;
  wire [31:0] icache_io_cpu_btb_update_bits_target;
  wire  icache_io_cpu_btb_update_bits_taken;
  wire  icache_io_cpu_btb_update_bits_isJump;
  wire  icache_io_cpu_btb_update_bits_isReturn;
  wire [31:0] icache_io_cpu_btb_update_bits_br_pc;
  wire  icache_io_cpu_bht_update_valid;
  wire  icache_io_cpu_bht_update_bits_prediction_valid;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_taken;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_mask;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_bridx;
  wire [31:0] icache_io_cpu_bht_update_bits_prediction_bits_target;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_entry;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_bht_history;
  wire [1:0] icache_io_cpu_bht_update_bits_prediction_bits_bht_value;
  wire [31:0] icache_io_cpu_bht_update_bits_pc;
  wire  icache_io_cpu_bht_update_bits_taken;
  wire  icache_io_cpu_bht_update_bits_mispredict;
  wire  icache_io_cpu_ras_update_valid;
  wire  icache_io_cpu_ras_update_bits_isCall;
  wire  icache_io_cpu_ras_update_bits_isReturn;
  wire [31:0] icache_io_cpu_ras_update_bits_returnAddr;
  wire  icache_io_cpu_ras_update_bits_prediction_valid;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_taken;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_mask;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_bridx;
  wire [31:0] icache_io_cpu_ras_update_bits_prediction_bits_target;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_entry;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_bht_history;
  wire [1:0] icache_io_cpu_ras_update_bits_prediction_bits_bht_value;
  wire  icache_io_cpu_flush_icache;
  wire  icache_io_cpu_flush_tlb;
  wire [31:0] icache_io_cpu_npc;
  wire  icache_io_ptw_req_ready;
  wire  icache_io_ptw_req_valid;
  wire [1:0] icache_io_ptw_req_bits_prv;
  wire  icache_io_ptw_req_bits_pum;
  wire  icache_io_ptw_req_bits_mxr;
  wire [19:0] icache_io_ptw_req_bits_addr;
  wire  icache_io_ptw_req_bits_store;
  wire  icache_io_ptw_req_bits_fetch;
  wire  icache_io_ptw_resp_valid;
  wire [15:0] icache_io_ptw_resp_bits_pte_reserved_for_hardware;
  wire [37:0] icache_io_ptw_resp_bits_pte_ppn;
  wire [1:0] icache_io_ptw_resp_bits_pte_reserved_for_software;
  wire  icache_io_ptw_resp_bits_pte_d;
  wire  icache_io_ptw_resp_bits_pte_a;
  wire  icache_io_ptw_resp_bits_pte_g;
  wire  icache_io_ptw_resp_bits_pte_u;
  wire  icache_io_ptw_resp_bits_pte_x;
  wire  icache_io_ptw_resp_bits_pte_w;
  wire  icache_io_ptw_resp_bits_pte_r;
  wire  icache_io_ptw_resp_bits_pte_v;
  wire [6:0] icache_io_ptw_ptbr_asid;
  wire [21:0] icache_io_ptw_ptbr_ppn;
  wire  icache_io_ptw_invalidate;
  wire  icache_io_ptw_status_debug;
  wire [1:0] icache_io_ptw_status_prv;
  wire  icache_io_ptw_status_sd;
  wire [30:0] icache_io_ptw_status_zero3;
  wire  icache_io_ptw_status_sd_rv32;
  wire [1:0] icache_io_ptw_status_zero2;
  wire [4:0] icache_io_ptw_status_vm;
  wire [3:0] icache_io_ptw_status_zero1;
  wire  icache_io_ptw_status_mxr;
  wire  icache_io_ptw_status_pum;
  wire  icache_io_ptw_status_mprv;
  wire [1:0] icache_io_ptw_status_xs;
  wire [1:0] icache_io_ptw_status_fs;
  wire [1:0] icache_io_ptw_status_mpp;
  wire [1:0] icache_io_ptw_status_hpp;
  wire  icache_io_ptw_status_spp;
  wire  icache_io_ptw_status_mpie;
  wire  icache_io_ptw_status_hpie;
  wire  icache_io_ptw_status_spie;
  wire  icache_io_ptw_status_upie;
  wire  icache_io_ptw_status_mie;
  wire  icache_io_ptw_status_hie;
  wire  icache_io_ptw_status_sie;
  wire  icache_io_ptw_status_uie;
  wire  icache_io_mem_acquire_ready;
  wire  icache_io_mem_acquire_valid;
  wire [25:0] icache_io_mem_acquire_bits_addr_block;
  wire  icache_io_mem_acquire_bits_client_xact_id;
  wire [2:0] icache_io_mem_acquire_bits_addr_beat;
  wire  icache_io_mem_acquire_bits_is_builtin_type;
  wire [2:0] icache_io_mem_acquire_bits_a_type;
  wire [11:0] icache_io_mem_acquire_bits_union;
  wire [63:0] icache_io_mem_acquire_bits_data;
  wire  icache_io_mem_grant_ready;
  wire  icache_io_mem_grant_valid;
  wire [2:0] icache_io_mem_grant_bits_addr_beat;
  wire  icache_io_mem_grant_bits_client_xact_id;
  wire [1:0] icache_io_mem_grant_bits_manager_xact_id;
  wire  icache_io_mem_grant_bits_is_builtin_type;
  wire [3:0] icache_io_mem_grant_bits_g_type;
  wire [63:0] icache_io_mem_grant_bits_data;
  wire  DCache_1_clk;
  wire  DCache_1_reset;
  wire  DCache_1_io_cpu_req_ready;
  wire  DCache_1_io_cpu_req_valid;
  wire [31:0] DCache_1_io_cpu_req_bits_addr;
  wire [8:0] DCache_1_io_cpu_req_bits_tag;
  wire [4:0] DCache_1_io_cpu_req_bits_cmd;
  wire [2:0] DCache_1_io_cpu_req_bits_typ;
  wire  DCache_1_io_cpu_req_bits_phys;
  wire [31:0] DCache_1_io_cpu_req_bits_data;
  wire  DCache_1_io_cpu_s1_kill;
  wire [31:0] DCache_1_io_cpu_s1_data;
  wire  DCache_1_io_cpu_s2_nack;
  wire  DCache_1_io_cpu_resp_valid;
  wire [31:0] DCache_1_io_cpu_resp_bits_addr;
  wire [8:0] DCache_1_io_cpu_resp_bits_tag;
  wire [4:0] DCache_1_io_cpu_resp_bits_cmd;
  wire [2:0] DCache_1_io_cpu_resp_bits_typ;
  wire [31:0] DCache_1_io_cpu_resp_bits_data;
  wire  DCache_1_io_cpu_resp_bits_replay;
  wire  DCache_1_io_cpu_resp_bits_has_data;
  wire [31:0] DCache_1_io_cpu_resp_bits_data_word_bypass;
  wire [31:0] DCache_1_io_cpu_resp_bits_store_data;
  wire  DCache_1_io_cpu_replay_next;
  wire  DCache_1_io_cpu_xcpt_ma_ld;
  wire  DCache_1_io_cpu_xcpt_ma_st;
  wire  DCache_1_io_cpu_xcpt_pf_ld;
  wire  DCache_1_io_cpu_xcpt_pf_st;
  wire  DCache_1_io_cpu_invalidate_lr;
  wire  DCache_1_io_cpu_ordered;
  wire  DCache_1_io_ptw_req_ready;
  wire  DCache_1_io_ptw_req_valid;
  wire [1:0] DCache_1_io_ptw_req_bits_prv;
  wire  DCache_1_io_ptw_req_bits_pum;
  wire  DCache_1_io_ptw_req_bits_mxr;
  wire [19:0] DCache_1_io_ptw_req_bits_addr;
  wire  DCache_1_io_ptw_req_bits_store;
  wire  DCache_1_io_ptw_req_bits_fetch;
  wire  DCache_1_io_ptw_resp_valid;
  wire [15:0] DCache_1_io_ptw_resp_bits_pte_reserved_for_hardware;
  wire [37:0] DCache_1_io_ptw_resp_bits_pte_ppn;
  wire [1:0] DCache_1_io_ptw_resp_bits_pte_reserved_for_software;
  wire  DCache_1_io_ptw_resp_bits_pte_d;
  wire  DCache_1_io_ptw_resp_bits_pte_a;
  wire  DCache_1_io_ptw_resp_bits_pte_g;
  wire  DCache_1_io_ptw_resp_bits_pte_u;
  wire  DCache_1_io_ptw_resp_bits_pte_x;
  wire  DCache_1_io_ptw_resp_bits_pte_w;
  wire  DCache_1_io_ptw_resp_bits_pte_r;
  wire  DCache_1_io_ptw_resp_bits_pte_v;
  wire [6:0] DCache_1_io_ptw_ptbr_asid;
  wire [21:0] DCache_1_io_ptw_ptbr_ppn;
  wire  DCache_1_io_ptw_invalidate;
  wire  DCache_1_io_ptw_status_debug;
  wire [1:0] DCache_1_io_ptw_status_prv;
  wire  DCache_1_io_ptw_status_sd;
  wire [30:0] DCache_1_io_ptw_status_zero3;
  wire  DCache_1_io_ptw_status_sd_rv32;
  wire [1:0] DCache_1_io_ptw_status_zero2;
  wire [4:0] DCache_1_io_ptw_status_vm;
  wire [3:0] DCache_1_io_ptw_status_zero1;
  wire  DCache_1_io_ptw_status_mxr;
  wire  DCache_1_io_ptw_status_pum;
  wire  DCache_1_io_ptw_status_mprv;
  wire [1:0] DCache_1_io_ptw_status_xs;
  wire [1:0] DCache_1_io_ptw_status_fs;
  wire [1:0] DCache_1_io_ptw_status_mpp;
  wire [1:0] DCache_1_io_ptw_status_hpp;
  wire  DCache_1_io_ptw_status_spp;
  wire  DCache_1_io_ptw_status_mpie;
  wire  DCache_1_io_ptw_status_hpie;
  wire  DCache_1_io_ptw_status_spie;
  wire  DCache_1_io_ptw_status_upie;
  wire  DCache_1_io_ptw_status_mie;
  wire  DCache_1_io_ptw_status_hie;
  wire  DCache_1_io_ptw_status_sie;
  wire  DCache_1_io_ptw_status_uie;
  wire  DCache_1_io_mem_acquire_ready;
  wire  DCache_1_io_mem_acquire_valid;
  wire [25:0] DCache_1_io_mem_acquire_bits_addr_block;
  wire  DCache_1_io_mem_acquire_bits_client_xact_id;
  wire [2:0] DCache_1_io_mem_acquire_bits_addr_beat;
  wire  DCache_1_io_mem_acquire_bits_is_builtin_type;
  wire [2:0] DCache_1_io_mem_acquire_bits_a_type;
  wire [11:0] DCache_1_io_mem_acquire_bits_union;
  wire [63:0] DCache_1_io_mem_acquire_bits_data;
  wire  DCache_1_io_mem_probe_ready;
  wire  DCache_1_io_mem_probe_valid;
  wire [25:0] DCache_1_io_mem_probe_bits_addr_block;
  wire [1:0] DCache_1_io_mem_probe_bits_p_type;
  wire  DCache_1_io_mem_release_ready;
  wire  DCache_1_io_mem_release_valid;
  wire [2:0] DCache_1_io_mem_release_bits_addr_beat;
  wire [25:0] DCache_1_io_mem_release_bits_addr_block;
  wire  DCache_1_io_mem_release_bits_client_xact_id;
  wire  DCache_1_io_mem_release_bits_voluntary;
  wire [2:0] DCache_1_io_mem_release_bits_r_type;
  wire [63:0] DCache_1_io_mem_release_bits_data;
  wire  DCache_1_io_mem_grant_ready;
  wire  DCache_1_io_mem_grant_valid;
  wire [2:0] DCache_1_io_mem_grant_bits_addr_beat;
  wire  DCache_1_io_mem_grant_bits_client_xact_id;
  wire [1:0] DCache_1_io_mem_grant_bits_manager_xact_id;
  wire  DCache_1_io_mem_grant_bits_is_builtin_type;
  wire [3:0] DCache_1_io_mem_grant_bits_g_type;
  wire [63:0] DCache_1_io_mem_grant_bits_data;
  wire  DCache_1_io_mem_grant_bits_manager_id;
  wire  DCache_1_io_mem_finish_ready;
  wire  DCache_1_io_mem_finish_valid;
  wire [1:0] DCache_1_io_mem_finish_bits_manager_xact_id;
  wire  DCache_1_io_mem_finish_bits_manager_id;
  wire  uncachedArb_clk;
  wire  uncachedArb_reset;
  wire  uncachedArb_io_in_0_acquire_ready;
  wire  uncachedArb_io_in_0_acquire_valid;
  wire [25:0] uncachedArb_io_in_0_acquire_bits_addr_block;
  wire  uncachedArb_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] uncachedArb_io_in_0_acquire_bits_addr_beat;
  wire  uncachedArb_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] uncachedArb_io_in_0_acquire_bits_a_type;
  wire [11:0] uncachedArb_io_in_0_acquire_bits_union;
  wire [63:0] uncachedArb_io_in_0_acquire_bits_data;
  wire  uncachedArb_io_in_0_grant_ready;
  wire  uncachedArb_io_in_0_grant_valid;
  wire [2:0] uncachedArb_io_in_0_grant_bits_addr_beat;
  wire  uncachedArb_io_in_0_grant_bits_client_xact_id;
  wire [1:0] uncachedArb_io_in_0_grant_bits_manager_xact_id;
  wire  uncachedArb_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] uncachedArb_io_in_0_grant_bits_g_type;
  wire [63:0] uncachedArb_io_in_0_grant_bits_data;
  wire  uncachedArb_io_out_acquire_ready;
  wire  uncachedArb_io_out_acquire_valid;
  wire [25:0] uncachedArb_io_out_acquire_bits_addr_block;
  wire  uncachedArb_io_out_acquire_bits_client_xact_id;
  wire [2:0] uncachedArb_io_out_acquire_bits_addr_beat;
  wire  uncachedArb_io_out_acquire_bits_is_builtin_type;
  wire [2:0] uncachedArb_io_out_acquire_bits_a_type;
  wire [11:0] uncachedArb_io_out_acquire_bits_union;
  wire [63:0] uncachedArb_io_out_acquire_bits_data;
  wire  uncachedArb_io_out_grant_ready;
  wire  uncachedArb_io_out_grant_valid;
  wire [2:0] uncachedArb_io_out_grant_bits_addr_beat;
  wire  uncachedArb_io_out_grant_bits_client_xact_id;
  wire [1:0] uncachedArb_io_out_grant_bits_manager_xact_id;
  wire  uncachedArb_io_out_grant_bits_is_builtin_type;
  wire [3:0] uncachedArb_io_out_grant_bits_g_type;
  wire [63:0] uncachedArb_io_out_grant_bits_data;
  wire  dcArb_clk;
  wire  dcArb_reset;
  wire  dcArb_io_requestor_0_req_ready;
  wire  dcArb_io_requestor_0_req_valid;
  wire [31:0] dcArb_io_requestor_0_req_bits_addr;
  wire [8:0] dcArb_io_requestor_0_req_bits_tag;
  wire [4:0] dcArb_io_requestor_0_req_bits_cmd;
  wire [2:0] dcArb_io_requestor_0_req_bits_typ;
  wire  dcArb_io_requestor_0_req_bits_phys;
  wire [31:0] dcArb_io_requestor_0_req_bits_data;
  wire  dcArb_io_requestor_0_s1_kill;
  wire [31:0] dcArb_io_requestor_0_s1_data;
  wire  dcArb_io_requestor_0_s2_nack;
  wire  dcArb_io_requestor_0_resp_valid;
  wire [31:0] dcArb_io_requestor_0_resp_bits_addr;
  wire [8:0] dcArb_io_requestor_0_resp_bits_tag;
  wire [4:0] dcArb_io_requestor_0_resp_bits_cmd;
  wire [2:0] dcArb_io_requestor_0_resp_bits_typ;
  wire [31:0] dcArb_io_requestor_0_resp_bits_data;
  wire  dcArb_io_requestor_0_resp_bits_replay;
  wire  dcArb_io_requestor_0_resp_bits_has_data;
  wire [31:0] dcArb_io_requestor_0_resp_bits_data_word_bypass;
  wire [31:0] dcArb_io_requestor_0_resp_bits_store_data;
  wire  dcArb_io_requestor_0_replay_next;
  wire  dcArb_io_requestor_0_xcpt_ma_ld;
  wire  dcArb_io_requestor_0_xcpt_ma_st;
  wire  dcArb_io_requestor_0_xcpt_pf_ld;
  wire  dcArb_io_requestor_0_xcpt_pf_st;
  wire  dcArb_io_requestor_0_invalidate_lr;
  wire  dcArb_io_requestor_0_ordered;
  wire  dcArb_io_mem_req_ready;
  wire  dcArb_io_mem_req_valid;
  wire [31:0] dcArb_io_mem_req_bits_addr;
  wire [8:0] dcArb_io_mem_req_bits_tag;
  wire [4:0] dcArb_io_mem_req_bits_cmd;
  wire [2:0] dcArb_io_mem_req_bits_typ;
  wire  dcArb_io_mem_req_bits_phys;
  wire [31:0] dcArb_io_mem_req_bits_data;
  wire  dcArb_io_mem_s1_kill;
  wire [31:0] dcArb_io_mem_s1_data;
  wire  dcArb_io_mem_s2_nack;
  wire  dcArb_io_mem_resp_valid;
  wire [31:0] dcArb_io_mem_resp_bits_addr;
  wire [8:0] dcArb_io_mem_resp_bits_tag;
  wire [4:0] dcArb_io_mem_resp_bits_cmd;
  wire [2:0] dcArb_io_mem_resp_bits_typ;
  wire [31:0] dcArb_io_mem_resp_bits_data;
  wire  dcArb_io_mem_resp_bits_replay;
  wire  dcArb_io_mem_resp_bits_has_data;
  wire [31:0] dcArb_io_mem_resp_bits_data_word_bypass;
  wire [31:0] dcArb_io_mem_resp_bits_store_data;
  wire  dcArb_io_mem_replay_next;
  wire  dcArb_io_mem_xcpt_ma_ld;
  wire  dcArb_io_mem_xcpt_ma_st;
  wire  dcArb_io_mem_xcpt_pf_ld;
  wire  dcArb_io_mem_xcpt_pf_st;
  wire  dcArb_io_mem_invalidate_lr;
  wire  dcArb_io_mem_ordered;
  reg  GEN_0;
  reg [31:0] GEN_160;
  reg [4:0] GEN_1;
  reg [31:0] GEN_161;
  reg [63:0] GEN_2;
  reg [63:0] GEN_162;
  reg [31:0] GEN_3;
  reg [31:0] GEN_163;
  reg  GEN_4;
  reg [31:0] GEN_164;
  reg  GEN_5;
  reg [31:0] GEN_165;
  reg  GEN_6;
  reg [31:0] GEN_166;
  reg [4:0] GEN_7;
  reg [31:0] GEN_167;
  reg  GEN_8;
  reg [31:0] GEN_168;
  reg  GEN_9;
  reg [31:0] GEN_169;
  reg  GEN_10;
  reg [31:0] GEN_170;
  reg  GEN_11;
  reg [31:0] GEN_171;
  reg  GEN_12;
  reg [31:0] GEN_172;
  reg  GEN_13;
  reg [31:0] GEN_173;
  reg  GEN_14;
  reg [31:0] GEN_174;
  reg  GEN_15;
  reg [31:0] GEN_175;
  reg  GEN_16;
  reg [31:0] GEN_176;
  reg  GEN_17;
  reg [31:0] GEN_177;
  reg  GEN_18;
  reg [31:0] GEN_178;
  reg  GEN_19;
  reg [31:0] GEN_179;
  reg  GEN_20;
  reg [31:0] GEN_180;
  reg  GEN_21;
  reg [31:0] GEN_181;
  reg  GEN_22;
  reg [31:0] GEN_182;
  reg  GEN_23;
  reg [31:0] GEN_183;
  reg  GEN_24;
  reg [31:0] GEN_184;
  reg  GEN_25;
  reg [31:0] GEN_185;
  reg [4:0] GEN_26;
  reg [31:0] GEN_186;
  reg  GEN_27;
  reg [31:0] GEN_187;
  reg  GEN_28;
  reg [31:0] GEN_188;
  reg [64:0] GEN_29;
  reg [95:0] GEN_189;
  reg [4:0] GEN_30;
  reg [31:0] GEN_190;
  reg  GEN_31;
  reg [31:0] GEN_191;
  reg  GEN_32;
  reg [31:0] GEN_192;
  reg [4:0] GEN_33;
  reg [31:0] GEN_193;
  reg [31:0] GEN_34;
  reg [31:0] GEN_194;
  reg  GEN_35;
  reg [31:0] GEN_195;
  reg [31:0] GEN_36;
  reg [31:0] GEN_196;
  reg [8:0] GEN_37;
  reg [31:0] GEN_197;
  reg [4:0] GEN_38;
  reg [31:0] GEN_198;
  reg [2:0] GEN_39;
  reg [31:0] GEN_199;
  reg  GEN_40;
  reg [31:0] GEN_200;
  reg [31:0] GEN_41;
  reg [31:0] GEN_201;
  reg  GEN_42;
  reg [31:0] GEN_202;
  reg [31:0] GEN_43;
  reg [31:0] GEN_203;
  reg  GEN_44;
  reg [31:0] GEN_204;
  reg  GEN_45;
  reg [31:0] GEN_205;
  reg  GEN_46;
  reg [31:0] GEN_206;
  reg  GEN_47;
  reg [31:0] GEN_207;
  reg [25:0] GEN_48;
  reg [31:0] GEN_208;
  reg  GEN_49;
  reg [31:0] GEN_209;
  reg [2:0] GEN_50;
  reg [31:0] GEN_210;
  reg  GEN_51;
  reg [31:0] GEN_211;
  reg [2:0] GEN_52;
  reg [31:0] GEN_212;
  reg [11:0] GEN_53;
  reg [31:0] GEN_213;
  reg [63:0] GEN_54;
  reg [63:0] GEN_214;
  reg  GEN_55;
  reg [31:0] GEN_215;
  reg  GEN_56;
  reg [31:0] GEN_216;
  reg [4:0] GEN_57;
  reg [31:0] GEN_217;
  reg  GEN_58;
  reg [31:0] GEN_218;
  reg  GEN_59;
  reg [31:0] GEN_219;
  reg  GEN_60;
  reg [31:0] GEN_220;
  reg  GEN_61;
  reg [31:0] GEN_221;
  reg  GEN_62;
  reg [31:0] GEN_222;
  reg  GEN_63;
  reg [31:0] GEN_223;
  reg  GEN_64;
  reg [31:0] GEN_224;
  reg  GEN_65;
  reg [31:0] GEN_225;
  reg  GEN_66;
  reg [31:0] GEN_226;
  reg  GEN_67;
  reg [31:0] GEN_227;
  reg  GEN_68;
  reg [31:0] GEN_228;
  reg  GEN_69;
  reg [31:0] GEN_229;
  reg  GEN_70;
  reg [31:0] GEN_230;
  reg  GEN_71;
  reg [31:0] GEN_231;
  reg  GEN_72;
  reg [31:0] GEN_232;
  reg  GEN_73;
  reg [31:0] GEN_233;
  reg [2:0] GEN_74;
  reg [31:0] GEN_234;
  reg [1:0] GEN_75;
  reg [31:0] GEN_235;
  reg [64:0] GEN_76;
  reg [95:0] GEN_236;
  reg [64:0] GEN_77;
  reg [95:0] GEN_237;
  reg [64:0] GEN_78;
  reg [95:0] GEN_238;
  reg  GEN_79;
  reg [31:0] GEN_239;
  reg  GEN_80;
  reg [31:0] GEN_240;
  reg  GEN_81;
  reg [31:0] GEN_241;
  reg [15:0] GEN_82;
  reg [31:0] GEN_242;
  reg [37:0] GEN_83;
  reg [63:0] GEN_243;
  reg [1:0] GEN_84;
  reg [31:0] GEN_244;
  reg  GEN_85;
  reg [31:0] GEN_245;
  reg  GEN_86;
  reg [31:0] GEN_246;
  reg  GEN_87;
  reg [31:0] GEN_247;
  reg  GEN_88;
  reg [31:0] GEN_248;
  reg  GEN_89;
  reg [31:0] GEN_249;
  reg  GEN_90;
  reg [31:0] GEN_250;
  reg  GEN_91;
  reg [31:0] GEN_251;
  reg  GEN_92;
  reg [31:0] GEN_252;
  reg [6:0] GEN_93;
  reg [31:0] GEN_253;
  reg [21:0] GEN_94;
  reg [31:0] GEN_254;
  reg  GEN_95;
  reg [31:0] GEN_255;
  reg  GEN_96;
  reg [31:0] GEN_256;
  reg [1:0] GEN_97;
  reg [31:0] GEN_257;
  reg  GEN_98;
  reg [31:0] GEN_258;
  reg [30:0] GEN_99;
  reg [31:0] GEN_259;
  reg  GEN_100;
  reg [31:0] GEN_260;
  reg [1:0] GEN_101;
  reg [31:0] GEN_261;
  reg [4:0] GEN_102;
  reg [31:0] GEN_262;
  reg [3:0] GEN_103;
  reg [31:0] GEN_263;
  reg  GEN_104;
  reg [31:0] GEN_264;
  reg  GEN_105;
  reg [31:0] GEN_265;
  reg  GEN_106;
  reg [31:0] GEN_266;
  reg [1:0] GEN_107;
  reg [31:0] GEN_267;
  reg [1:0] GEN_108;
  reg [31:0] GEN_268;
  reg [1:0] GEN_109;
  reg [31:0] GEN_269;
  reg [1:0] GEN_110;
  reg [31:0] GEN_270;
  reg  GEN_111;
  reg [31:0] GEN_271;
  reg  GEN_112;
  reg [31:0] GEN_272;
  reg  GEN_113;
  reg [31:0] GEN_273;
  reg  GEN_114;
  reg [31:0] GEN_274;
  reg  GEN_115;
  reg [31:0] GEN_275;
  reg  GEN_116;
  reg [31:0] GEN_276;
  reg  GEN_117;
  reg [31:0] GEN_277;
  reg  GEN_118;
  reg [31:0] GEN_278;
  reg  GEN_119;
  reg [31:0] GEN_279;
  reg  GEN_120;
  reg [31:0] GEN_280;
  reg  GEN_121;
  reg [31:0] GEN_281;
  reg [15:0] GEN_122;
  reg [31:0] GEN_282;
  reg [37:0] GEN_123;
  reg [63:0] GEN_283;
  reg [1:0] GEN_124;
  reg [31:0] GEN_284;
  reg  GEN_125;
  reg [31:0] GEN_285;
  reg  GEN_126;
  reg [31:0] GEN_286;
  reg  GEN_127;
  reg [31:0] GEN_287;
  reg  GEN_128;
  reg [31:0] GEN_288;
  reg  GEN_129;
  reg [31:0] GEN_289;
  reg  GEN_130;
  reg [31:0] GEN_290;
  reg  GEN_131;
  reg [31:0] GEN_291;
  reg  GEN_132;
  reg [31:0] GEN_292;
  reg [6:0] GEN_133;
  reg [31:0] GEN_293;
  reg [21:0] GEN_134;
  reg [31:0] GEN_294;
  reg  GEN_135;
  reg [31:0] GEN_295;
  reg  GEN_136;
  reg [31:0] GEN_296;
  reg [1:0] GEN_137;
  reg [31:0] GEN_297;
  reg  GEN_138;
  reg [31:0] GEN_298;
  reg [30:0] GEN_139;
  reg [31:0] GEN_299;
  reg  GEN_140;
  reg [31:0] GEN_300;
  reg [1:0] GEN_141;
  reg [31:0] GEN_301;
  reg [4:0] GEN_142;
  reg [31:0] GEN_302;
  reg [3:0] GEN_143;
  reg [31:0] GEN_303;
  reg  GEN_144;
  reg [31:0] GEN_304;
  reg  GEN_145;
  reg [31:0] GEN_305;
  reg  GEN_146;
  reg [31:0] GEN_306;
  reg [1:0] GEN_147;
  reg [31:0] GEN_307;
  reg [1:0] GEN_148;
  reg [31:0] GEN_308;
  reg [1:0] GEN_149;
  reg [31:0] GEN_309;
  reg [1:0] GEN_150;
  reg [31:0] GEN_310;
  reg  GEN_151;
  reg [31:0] GEN_311;
  reg  GEN_152;
  reg [31:0] GEN_312;
  reg  GEN_153;
  reg [31:0] GEN_313;
  reg  GEN_154;
  reg [31:0] GEN_314;
  reg  GEN_155;
  reg [31:0] GEN_315;
  reg  GEN_156;
  reg [31:0] GEN_316;
  reg  GEN_157;
  reg [31:0] GEN_317;
  reg  GEN_158;
  reg [31:0] GEN_318;
  reg  GEN_159;
  reg [31:0] GEN_319;
  Rocket core (
    .clk(core_clk),
    .reset(core_reset),
    .io_prci_reset(core_io_prci_reset),
    .io_prci_id(core_io_prci_id),
    .io_prci_interrupts_meip(core_io_prci_interrupts_meip),
    .io_prci_interrupts_seip(core_io_prci_interrupts_seip),
    .io_prci_interrupts_debug(core_io_prci_interrupts_debug),
    .io_prci_interrupts_mtip(core_io_prci_interrupts_mtip),
    .io_prci_interrupts_msip(core_io_prci_interrupts_msip),
    .io_imem_req_valid(core_io_imem_req_valid),
    .io_imem_req_bits_pc(core_io_imem_req_bits_pc),
    .io_imem_req_bits_speculative(core_io_imem_req_bits_speculative),
    .io_imem_resp_ready(core_io_imem_resp_ready),
    .io_imem_resp_valid(core_io_imem_resp_valid),
    .io_imem_resp_bits_pc(core_io_imem_resp_bits_pc),
    .io_imem_resp_bits_data_0(core_io_imem_resp_bits_data_0),
    .io_imem_resp_bits_mask(core_io_imem_resp_bits_mask),
    .io_imem_resp_bits_xcpt_if(core_io_imem_resp_bits_xcpt_if),
    .io_imem_resp_bits_replay(core_io_imem_resp_bits_replay),
    .io_imem_btb_resp_valid(core_io_imem_btb_resp_valid),
    .io_imem_btb_resp_bits_taken(core_io_imem_btb_resp_bits_taken),
    .io_imem_btb_resp_bits_mask(core_io_imem_btb_resp_bits_mask),
    .io_imem_btb_resp_bits_bridx(core_io_imem_btb_resp_bits_bridx),
    .io_imem_btb_resp_bits_target(core_io_imem_btb_resp_bits_target),
    .io_imem_btb_resp_bits_entry(core_io_imem_btb_resp_bits_entry),
    .io_imem_btb_resp_bits_bht_history(core_io_imem_btb_resp_bits_bht_history),
    .io_imem_btb_resp_bits_bht_value(core_io_imem_btb_resp_bits_bht_value),
    .io_imem_btb_update_valid(core_io_imem_btb_update_valid),
    .io_imem_btb_update_bits_prediction_valid(core_io_imem_btb_update_bits_prediction_valid),
    .io_imem_btb_update_bits_prediction_bits_taken(core_io_imem_btb_update_bits_prediction_bits_taken),
    .io_imem_btb_update_bits_prediction_bits_mask(core_io_imem_btb_update_bits_prediction_bits_mask),
    .io_imem_btb_update_bits_prediction_bits_bridx(core_io_imem_btb_update_bits_prediction_bits_bridx),
    .io_imem_btb_update_bits_prediction_bits_target(core_io_imem_btb_update_bits_prediction_bits_target),
    .io_imem_btb_update_bits_prediction_bits_entry(core_io_imem_btb_update_bits_prediction_bits_entry),
    .io_imem_btb_update_bits_prediction_bits_bht_history(core_io_imem_btb_update_bits_prediction_bits_bht_history),
    .io_imem_btb_update_bits_prediction_bits_bht_value(core_io_imem_btb_update_bits_prediction_bits_bht_value),
    .io_imem_btb_update_bits_pc(core_io_imem_btb_update_bits_pc),
    .io_imem_btb_update_bits_target(core_io_imem_btb_update_bits_target),
    .io_imem_btb_update_bits_taken(core_io_imem_btb_update_bits_taken),
    .io_imem_btb_update_bits_isJump(core_io_imem_btb_update_bits_isJump),
    .io_imem_btb_update_bits_isReturn(core_io_imem_btb_update_bits_isReturn),
    .io_imem_btb_update_bits_br_pc(core_io_imem_btb_update_bits_br_pc),
    .io_imem_bht_update_valid(core_io_imem_bht_update_valid),
    .io_imem_bht_update_bits_prediction_valid(core_io_imem_bht_update_bits_prediction_valid),
    .io_imem_bht_update_bits_prediction_bits_taken(core_io_imem_bht_update_bits_prediction_bits_taken),
    .io_imem_bht_update_bits_prediction_bits_mask(core_io_imem_bht_update_bits_prediction_bits_mask),
    .io_imem_bht_update_bits_prediction_bits_bridx(core_io_imem_bht_update_bits_prediction_bits_bridx),
    .io_imem_bht_update_bits_prediction_bits_target(core_io_imem_bht_update_bits_prediction_bits_target),
    .io_imem_bht_update_bits_prediction_bits_entry(core_io_imem_bht_update_bits_prediction_bits_entry),
    .io_imem_bht_update_bits_prediction_bits_bht_history(core_io_imem_bht_update_bits_prediction_bits_bht_history),
    .io_imem_bht_update_bits_prediction_bits_bht_value(core_io_imem_bht_update_bits_prediction_bits_bht_value),
    .io_imem_bht_update_bits_pc(core_io_imem_bht_update_bits_pc),
    .io_imem_bht_update_bits_taken(core_io_imem_bht_update_bits_taken),
    .io_imem_bht_update_bits_mispredict(core_io_imem_bht_update_bits_mispredict),
    .io_imem_ras_update_valid(core_io_imem_ras_update_valid),
    .io_imem_ras_update_bits_isCall(core_io_imem_ras_update_bits_isCall),
    .io_imem_ras_update_bits_isReturn(core_io_imem_ras_update_bits_isReturn),
    .io_imem_ras_update_bits_returnAddr(core_io_imem_ras_update_bits_returnAddr),
    .io_imem_ras_update_bits_prediction_valid(core_io_imem_ras_update_bits_prediction_valid),
    .io_imem_ras_update_bits_prediction_bits_taken(core_io_imem_ras_update_bits_prediction_bits_taken),
    .io_imem_ras_update_bits_prediction_bits_mask(core_io_imem_ras_update_bits_prediction_bits_mask),
    .io_imem_ras_update_bits_prediction_bits_bridx(core_io_imem_ras_update_bits_prediction_bits_bridx),
    .io_imem_ras_update_bits_prediction_bits_target(core_io_imem_ras_update_bits_prediction_bits_target),
    .io_imem_ras_update_bits_prediction_bits_entry(core_io_imem_ras_update_bits_prediction_bits_entry),
    .io_imem_ras_update_bits_prediction_bits_bht_history(core_io_imem_ras_update_bits_prediction_bits_bht_history),
    .io_imem_ras_update_bits_prediction_bits_bht_value(core_io_imem_ras_update_bits_prediction_bits_bht_value),
    .io_imem_flush_icache(core_io_imem_flush_icache),
    .io_imem_flush_tlb(core_io_imem_flush_tlb),
    .io_imem_npc(core_io_imem_npc),
    .io_dmem_req_ready(core_io_dmem_req_ready),
    .io_dmem_req_valid(core_io_dmem_req_valid),
    .io_dmem_req_bits_addr(core_io_dmem_req_bits_addr),
    .io_dmem_req_bits_tag(core_io_dmem_req_bits_tag),
    .io_dmem_req_bits_cmd(core_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_typ(core_io_dmem_req_bits_typ),
    .io_dmem_req_bits_phys(core_io_dmem_req_bits_phys),
    .io_dmem_req_bits_data(core_io_dmem_req_bits_data),
    .io_dmem_s1_kill(core_io_dmem_s1_kill),
    .io_dmem_s1_data(core_io_dmem_s1_data),
    .io_dmem_s2_nack(core_io_dmem_s2_nack),
    .io_dmem_resp_valid(core_io_dmem_resp_valid),
    .io_dmem_resp_bits_addr(core_io_dmem_resp_bits_addr),
    .io_dmem_resp_bits_tag(core_io_dmem_resp_bits_tag),
    .io_dmem_resp_bits_cmd(core_io_dmem_resp_bits_cmd),
    .io_dmem_resp_bits_typ(core_io_dmem_resp_bits_typ),
    .io_dmem_resp_bits_data(core_io_dmem_resp_bits_data),
    .io_dmem_resp_bits_replay(core_io_dmem_resp_bits_replay),
    .io_dmem_resp_bits_has_data(core_io_dmem_resp_bits_has_data),
    .io_dmem_resp_bits_data_word_bypass(core_io_dmem_resp_bits_data_word_bypass),
    .io_dmem_resp_bits_store_data(core_io_dmem_resp_bits_store_data),
    .io_dmem_replay_next(core_io_dmem_replay_next),
    .io_dmem_xcpt_ma_ld(core_io_dmem_xcpt_ma_ld),
    .io_dmem_xcpt_ma_st(core_io_dmem_xcpt_ma_st),
    .io_dmem_xcpt_pf_ld(core_io_dmem_xcpt_pf_ld),
    .io_dmem_xcpt_pf_st(core_io_dmem_xcpt_pf_st),
    .io_dmem_invalidate_lr(core_io_dmem_invalidate_lr),
    .io_dmem_ordered(core_io_dmem_ordered),
    .io_ptw_ptbr_asid(core_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(core_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(core_io_ptw_invalidate),
    .io_ptw_status_debug(core_io_ptw_status_debug),
    .io_ptw_status_prv(core_io_ptw_status_prv),
    .io_ptw_status_sd(core_io_ptw_status_sd),
    .io_ptw_status_zero3(core_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(core_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(core_io_ptw_status_zero2),
    .io_ptw_status_vm(core_io_ptw_status_vm),
    .io_ptw_status_zero1(core_io_ptw_status_zero1),
    .io_ptw_status_mxr(core_io_ptw_status_mxr),
    .io_ptw_status_pum(core_io_ptw_status_pum),
    .io_ptw_status_mprv(core_io_ptw_status_mprv),
    .io_ptw_status_xs(core_io_ptw_status_xs),
    .io_ptw_status_fs(core_io_ptw_status_fs),
    .io_ptw_status_mpp(core_io_ptw_status_mpp),
    .io_ptw_status_hpp(core_io_ptw_status_hpp),
    .io_ptw_status_spp(core_io_ptw_status_spp),
    .io_ptw_status_mpie(core_io_ptw_status_mpie),
    .io_ptw_status_hpie(core_io_ptw_status_hpie),
    .io_ptw_status_spie(core_io_ptw_status_spie),
    .io_ptw_status_upie(core_io_ptw_status_upie),
    .io_ptw_status_mie(core_io_ptw_status_mie),
    .io_ptw_status_hie(core_io_ptw_status_hie),
    .io_ptw_status_sie(core_io_ptw_status_sie),
    .io_ptw_status_uie(core_io_ptw_status_uie),
    .io_fpu_inst(core_io_fpu_inst),
    .io_fpu_fromint_data(core_io_fpu_fromint_data),
    .io_fpu_fcsr_rm(core_io_fpu_fcsr_rm),
    .io_fpu_fcsr_flags_valid(core_io_fpu_fcsr_flags_valid),
    .io_fpu_fcsr_flags_bits(core_io_fpu_fcsr_flags_bits),
    .io_fpu_store_data(core_io_fpu_store_data),
    .io_fpu_toint_data(core_io_fpu_toint_data),
    .io_fpu_dmem_resp_val(core_io_fpu_dmem_resp_val),
    .io_fpu_dmem_resp_type(core_io_fpu_dmem_resp_type),
    .io_fpu_dmem_resp_tag(core_io_fpu_dmem_resp_tag),
    .io_fpu_dmem_resp_data(core_io_fpu_dmem_resp_data),
    .io_fpu_valid(core_io_fpu_valid),
    .io_fpu_fcsr_rdy(core_io_fpu_fcsr_rdy),
    .io_fpu_nack_mem(core_io_fpu_nack_mem),
    .io_fpu_illegal_rm(core_io_fpu_illegal_rm),
    .io_fpu_killx(core_io_fpu_killx),
    .io_fpu_killm(core_io_fpu_killm),
    .io_fpu_dec_cmd(core_io_fpu_dec_cmd),
    .io_fpu_dec_ldst(core_io_fpu_dec_ldst),
    .io_fpu_dec_wen(core_io_fpu_dec_wen),
    .io_fpu_dec_ren1(core_io_fpu_dec_ren1),
    .io_fpu_dec_ren2(core_io_fpu_dec_ren2),
    .io_fpu_dec_ren3(core_io_fpu_dec_ren3),
    .io_fpu_dec_swap12(core_io_fpu_dec_swap12),
    .io_fpu_dec_swap23(core_io_fpu_dec_swap23),
    .io_fpu_dec_single(core_io_fpu_dec_single),
    .io_fpu_dec_fromint(core_io_fpu_dec_fromint),
    .io_fpu_dec_toint(core_io_fpu_dec_toint),
    .io_fpu_dec_fastpipe(core_io_fpu_dec_fastpipe),
    .io_fpu_dec_fma(core_io_fpu_dec_fma),
    .io_fpu_dec_div(core_io_fpu_dec_div),
    .io_fpu_dec_sqrt(core_io_fpu_dec_sqrt),
    .io_fpu_dec_round(core_io_fpu_dec_round),
    .io_fpu_dec_wflags(core_io_fpu_dec_wflags),
    .io_fpu_sboard_set(core_io_fpu_sboard_set),
    .io_fpu_sboard_clr(core_io_fpu_sboard_clr),
    .io_fpu_sboard_clra(core_io_fpu_sboard_clra),
    .io_fpu_cp_req_ready(core_io_fpu_cp_req_ready),
    .io_fpu_cp_req_valid(core_io_fpu_cp_req_valid),
    .io_fpu_cp_req_bits_cmd(core_io_fpu_cp_req_bits_cmd),
    .io_fpu_cp_req_bits_ldst(core_io_fpu_cp_req_bits_ldst),
    .io_fpu_cp_req_bits_wen(core_io_fpu_cp_req_bits_wen),
    .io_fpu_cp_req_bits_ren1(core_io_fpu_cp_req_bits_ren1),
    .io_fpu_cp_req_bits_ren2(core_io_fpu_cp_req_bits_ren2),
    .io_fpu_cp_req_bits_ren3(core_io_fpu_cp_req_bits_ren3),
    .io_fpu_cp_req_bits_swap12(core_io_fpu_cp_req_bits_swap12),
    .io_fpu_cp_req_bits_swap23(core_io_fpu_cp_req_bits_swap23),
    .io_fpu_cp_req_bits_single(core_io_fpu_cp_req_bits_single),
    .io_fpu_cp_req_bits_fromint(core_io_fpu_cp_req_bits_fromint),
    .io_fpu_cp_req_bits_toint(core_io_fpu_cp_req_bits_toint),
    .io_fpu_cp_req_bits_fastpipe(core_io_fpu_cp_req_bits_fastpipe),
    .io_fpu_cp_req_bits_fma(core_io_fpu_cp_req_bits_fma),
    .io_fpu_cp_req_bits_div(core_io_fpu_cp_req_bits_div),
    .io_fpu_cp_req_bits_sqrt(core_io_fpu_cp_req_bits_sqrt),
    .io_fpu_cp_req_bits_round(core_io_fpu_cp_req_bits_round),
    .io_fpu_cp_req_bits_wflags(core_io_fpu_cp_req_bits_wflags),
    .io_fpu_cp_req_bits_rm(core_io_fpu_cp_req_bits_rm),
    .io_fpu_cp_req_bits_typ(core_io_fpu_cp_req_bits_typ),
    .io_fpu_cp_req_bits_in1(core_io_fpu_cp_req_bits_in1),
    .io_fpu_cp_req_bits_in2(core_io_fpu_cp_req_bits_in2),
    .io_fpu_cp_req_bits_in3(core_io_fpu_cp_req_bits_in3),
    .io_fpu_cp_resp_ready(core_io_fpu_cp_resp_ready),
    .io_fpu_cp_resp_valid(core_io_fpu_cp_resp_valid),
    .io_fpu_cp_resp_bits_data(core_io_fpu_cp_resp_bits_data),
    .io_fpu_cp_resp_bits_exc(core_io_fpu_cp_resp_bits_exc),
    .io_rocc_cmd_ready(core_io_rocc_cmd_ready),
    .io_rocc_cmd_valid(core_io_rocc_cmd_valid),
    .io_rocc_cmd_bits_inst_funct(core_io_rocc_cmd_bits_inst_funct),
    .io_rocc_cmd_bits_inst_rs2(core_io_rocc_cmd_bits_inst_rs2),
    .io_rocc_cmd_bits_inst_rs1(core_io_rocc_cmd_bits_inst_rs1),
    .io_rocc_cmd_bits_inst_xd(core_io_rocc_cmd_bits_inst_xd),
    .io_rocc_cmd_bits_inst_xs1(core_io_rocc_cmd_bits_inst_xs1),
    .io_rocc_cmd_bits_inst_xs2(core_io_rocc_cmd_bits_inst_xs2),
    .io_rocc_cmd_bits_inst_rd(core_io_rocc_cmd_bits_inst_rd),
    .io_rocc_cmd_bits_inst_opcode(core_io_rocc_cmd_bits_inst_opcode),
    .io_rocc_cmd_bits_rs1(core_io_rocc_cmd_bits_rs1),
    .io_rocc_cmd_bits_rs2(core_io_rocc_cmd_bits_rs2),
    .io_rocc_cmd_bits_status_debug(core_io_rocc_cmd_bits_status_debug),
    .io_rocc_cmd_bits_status_prv(core_io_rocc_cmd_bits_status_prv),
    .io_rocc_cmd_bits_status_sd(core_io_rocc_cmd_bits_status_sd),
    .io_rocc_cmd_bits_status_zero3(core_io_rocc_cmd_bits_status_zero3),
    .io_rocc_cmd_bits_status_sd_rv32(core_io_rocc_cmd_bits_status_sd_rv32),
    .io_rocc_cmd_bits_status_zero2(core_io_rocc_cmd_bits_status_zero2),
    .io_rocc_cmd_bits_status_vm(core_io_rocc_cmd_bits_status_vm),
    .io_rocc_cmd_bits_status_zero1(core_io_rocc_cmd_bits_status_zero1),
    .io_rocc_cmd_bits_status_mxr(core_io_rocc_cmd_bits_status_mxr),
    .io_rocc_cmd_bits_status_pum(core_io_rocc_cmd_bits_status_pum),
    .io_rocc_cmd_bits_status_mprv(core_io_rocc_cmd_bits_status_mprv),
    .io_rocc_cmd_bits_status_xs(core_io_rocc_cmd_bits_status_xs),
    .io_rocc_cmd_bits_status_fs(core_io_rocc_cmd_bits_status_fs),
    .io_rocc_cmd_bits_status_mpp(core_io_rocc_cmd_bits_status_mpp),
    .io_rocc_cmd_bits_status_hpp(core_io_rocc_cmd_bits_status_hpp),
    .io_rocc_cmd_bits_status_spp(core_io_rocc_cmd_bits_status_spp),
    .io_rocc_cmd_bits_status_mpie(core_io_rocc_cmd_bits_status_mpie),
    .io_rocc_cmd_bits_status_hpie(core_io_rocc_cmd_bits_status_hpie),
    .io_rocc_cmd_bits_status_spie(core_io_rocc_cmd_bits_status_spie),
    .io_rocc_cmd_bits_status_upie(core_io_rocc_cmd_bits_status_upie),
    .io_rocc_cmd_bits_status_mie(core_io_rocc_cmd_bits_status_mie),
    .io_rocc_cmd_bits_status_hie(core_io_rocc_cmd_bits_status_hie),
    .io_rocc_cmd_bits_status_sie(core_io_rocc_cmd_bits_status_sie),
    .io_rocc_cmd_bits_status_uie(core_io_rocc_cmd_bits_status_uie),
    .io_rocc_resp_ready(core_io_rocc_resp_ready),
    .io_rocc_resp_valid(core_io_rocc_resp_valid),
    .io_rocc_resp_bits_rd(core_io_rocc_resp_bits_rd),
    .io_rocc_resp_bits_data(core_io_rocc_resp_bits_data),
    .io_rocc_mem_req_ready(core_io_rocc_mem_req_ready),
    .io_rocc_mem_req_valid(core_io_rocc_mem_req_valid),
    .io_rocc_mem_req_bits_addr(core_io_rocc_mem_req_bits_addr),
    .io_rocc_mem_req_bits_tag(core_io_rocc_mem_req_bits_tag),
    .io_rocc_mem_req_bits_cmd(core_io_rocc_mem_req_bits_cmd),
    .io_rocc_mem_req_bits_typ(core_io_rocc_mem_req_bits_typ),
    .io_rocc_mem_req_bits_phys(core_io_rocc_mem_req_bits_phys),
    .io_rocc_mem_req_bits_data(core_io_rocc_mem_req_bits_data),
    .io_rocc_mem_s1_kill(core_io_rocc_mem_s1_kill),
    .io_rocc_mem_s1_data(core_io_rocc_mem_s1_data),
    .io_rocc_mem_s2_nack(core_io_rocc_mem_s2_nack),
    .io_rocc_mem_resp_valid(core_io_rocc_mem_resp_valid),
    .io_rocc_mem_resp_bits_addr(core_io_rocc_mem_resp_bits_addr),
    .io_rocc_mem_resp_bits_tag(core_io_rocc_mem_resp_bits_tag),
    .io_rocc_mem_resp_bits_cmd(core_io_rocc_mem_resp_bits_cmd),
    .io_rocc_mem_resp_bits_typ(core_io_rocc_mem_resp_bits_typ),
    .io_rocc_mem_resp_bits_data(core_io_rocc_mem_resp_bits_data),
    .io_rocc_mem_resp_bits_replay(core_io_rocc_mem_resp_bits_replay),
    .io_rocc_mem_resp_bits_has_data(core_io_rocc_mem_resp_bits_has_data),
    .io_rocc_mem_resp_bits_data_word_bypass(core_io_rocc_mem_resp_bits_data_word_bypass),
    .io_rocc_mem_resp_bits_store_data(core_io_rocc_mem_resp_bits_store_data),
    .io_rocc_mem_replay_next(core_io_rocc_mem_replay_next),
    .io_rocc_mem_xcpt_ma_ld(core_io_rocc_mem_xcpt_ma_ld),
    .io_rocc_mem_xcpt_ma_st(core_io_rocc_mem_xcpt_ma_st),
    .io_rocc_mem_xcpt_pf_ld(core_io_rocc_mem_xcpt_pf_ld),
    .io_rocc_mem_xcpt_pf_st(core_io_rocc_mem_xcpt_pf_st),
    .io_rocc_mem_invalidate_lr(core_io_rocc_mem_invalidate_lr),
    .io_rocc_mem_ordered(core_io_rocc_mem_ordered),
    .io_rocc_busy(core_io_rocc_busy),
    .io_rocc_interrupt(core_io_rocc_interrupt),
    .io_rocc_autl_acquire_ready(core_io_rocc_autl_acquire_ready),
    .io_rocc_autl_acquire_valid(core_io_rocc_autl_acquire_valid),
    .io_rocc_autl_acquire_bits_addr_block(core_io_rocc_autl_acquire_bits_addr_block),
    .io_rocc_autl_acquire_bits_client_xact_id(core_io_rocc_autl_acquire_bits_client_xact_id),
    .io_rocc_autl_acquire_bits_addr_beat(core_io_rocc_autl_acquire_bits_addr_beat),
    .io_rocc_autl_acquire_bits_is_builtin_type(core_io_rocc_autl_acquire_bits_is_builtin_type),
    .io_rocc_autl_acquire_bits_a_type(core_io_rocc_autl_acquire_bits_a_type),
    .io_rocc_autl_acquire_bits_union(core_io_rocc_autl_acquire_bits_union),
    .io_rocc_autl_acquire_bits_data(core_io_rocc_autl_acquire_bits_data),
    .io_rocc_autl_grant_ready(core_io_rocc_autl_grant_ready),
    .io_rocc_autl_grant_valid(core_io_rocc_autl_grant_valid),
    .io_rocc_autl_grant_bits_addr_beat(core_io_rocc_autl_grant_bits_addr_beat),
    .io_rocc_autl_grant_bits_client_xact_id(core_io_rocc_autl_grant_bits_client_xact_id),
    .io_rocc_autl_grant_bits_manager_xact_id(core_io_rocc_autl_grant_bits_manager_xact_id),
    .io_rocc_autl_grant_bits_is_builtin_type(core_io_rocc_autl_grant_bits_is_builtin_type),
    .io_rocc_autl_grant_bits_g_type(core_io_rocc_autl_grant_bits_g_type),
    .io_rocc_autl_grant_bits_data(core_io_rocc_autl_grant_bits_data),
    .io_rocc_fpu_req_ready(core_io_rocc_fpu_req_ready),
    .io_rocc_fpu_req_valid(core_io_rocc_fpu_req_valid),
    .io_rocc_fpu_req_bits_cmd(core_io_rocc_fpu_req_bits_cmd),
    .io_rocc_fpu_req_bits_ldst(core_io_rocc_fpu_req_bits_ldst),
    .io_rocc_fpu_req_bits_wen(core_io_rocc_fpu_req_bits_wen),
    .io_rocc_fpu_req_bits_ren1(core_io_rocc_fpu_req_bits_ren1),
    .io_rocc_fpu_req_bits_ren2(core_io_rocc_fpu_req_bits_ren2),
    .io_rocc_fpu_req_bits_ren3(core_io_rocc_fpu_req_bits_ren3),
    .io_rocc_fpu_req_bits_swap12(core_io_rocc_fpu_req_bits_swap12),
    .io_rocc_fpu_req_bits_swap23(core_io_rocc_fpu_req_bits_swap23),
    .io_rocc_fpu_req_bits_single(core_io_rocc_fpu_req_bits_single),
    .io_rocc_fpu_req_bits_fromint(core_io_rocc_fpu_req_bits_fromint),
    .io_rocc_fpu_req_bits_toint(core_io_rocc_fpu_req_bits_toint),
    .io_rocc_fpu_req_bits_fastpipe(core_io_rocc_fpu_req_bits_fastpipe),
    .io_rocc_fpu_req_bits_fma(core_io_rocc_fpu_req_bits_fma),
    .io_rocc_fpu_req_bits_div(core_io_rocc_fpu_req_bits_div),
    .io_rocc_fpu_req_bits_sqrt(core_io_rocc_fpu_req_bits_sqrt),
    .io_rocc_fpu_req_bits_round(core_io_rocc_fpu_req_bits_round),
    .io_rocc_fpu_req_bits_wflags(core_io_rocc_fpu_req_bits_wflags),
    .io_rocc_fpu_req_bits_rm(core_io_rocc_fpu_req_bits_rm),
    .io_rocc_fpu_req_bits_typ(core_io_rocc_fpu_req_bits_typ),
    .io_rocc_fpu_req_bits_in1(core_io_rocc_fpu_req_bits_in1),
    .io_rocc_fpu_req_bits_in2(core_io_rocc_fpu_req_bits_in2),
    .io_rocc_fpu_req_bits_in3(core_io_rocc_fpu_req_bits_in3),
    .io_rocc_fpu_resp_ready(core_io_rocc_fpu_resp_ready),
    .io_rocc_fpu_resp_valid(core_io_rocc_fpu_resp_valid),
    .io_rocc_fpu_resp_bits_data(core_io_rocc_fpu_resp_bits_data),
    .io_rocc_fpu_resp_bits_exc(core_io_rocc_fpu_resp_bits_exc),
    .io_rocc_exception(core_io_rocc_exception),
    .io_rocc_csr_waddr(core_io_rocc_csr_waddr),
    .io_rocc_csr_wdata(core_io_rocc_csr_wdata),
    .io_rocc_csr_wen(core_io_rocc_csr_wen),
    .io_rocc_host_id(core_io_rocc_host_id)
  );
  
  //<CJ> RESET_VECTOR_ADDR
   defparam icache.RESET_VECTOR_ADDR = RESET_VECTOR_ADDR;
  
  Frontend icache (
    .clk(icache_clk),
    .reset(icache_reset),
    .io_cpu_req_valid(icache_io_cpu_req_valid),
    .io_cpu_req_bits_pc(icache_io_cpu_req_bits_pc),
    .io_cpu_req_bits_speculative(icache_io_cpu_req_bits_speculative),
    .io_cpu_resp_ready(icache_io_cpu_resp_ready),
    .io_cpu_resp_valid(icache_io_cpu_resp_valid),
    .io_cpu_resp_bits_pc(icache_io_cpu_resp_bits_pc),
    .io_cpu_resp_bits_data_0(icache_io_cpu_resp_bits_data_0),
    .io_cpu_resp_bits_mask(icache_io_cpu_resp_bits_mask),
    .io_cpu_resp_bits_xcpt_if(icache_io_cpu_resp_bits_xcpt_if),
    .io_cpu_resp_bits_replay(icache_io_cpu_resp_bits_replay),
    .io_cpu_btb_resp_valid(icache_io_cpu_btb_resp_valid),
    .io_cpu_btb_resp_bits_taken(icache_io_cpu_btb_resp_bits_taken),
    .io_cpu_btb_resp_bits_mask(icache_io_cpu_btb_resp_bits_mask),
    .io_cpu_btb_resp_bits_bridx(icache_io_cpu_btb_resp_bits_bridx),
    .io_cpu_btb_resp_bits_target(icache_io_cpu_btb_resp_bits_target),
    .io_cpu_btb_resp_bits_entry(icache_io_cpu_btb_resp_bits_entry),
    .io_cpu_btb_resp_bits_bht_history(icache_io_cpu_btb_resp_bits_bht_history),
    .io_cpu_btb_resp_bits_bht_value(icache_io_cpu_btb_resp_bits_bht_value),
    .io_cpu_btb_update_valid(icache_io_cpu_btb_update_valid),
    .io_cpu_btb_update_bits_prediction_valid(icache_io_cpu_btb_update_bits_prediction_valid),
    .io_cpu_btb_update_bits_prediction_bits_taken(icache_io_cpu_btb_update_bits_prediction_bits_taken),
    .io_cpu_btb_update_bits_prediction_bits_mask(icache_io_cpu_btb_update_bits_prediction_bits_mask),
    .io_cpu_btb_update_bits_prediction_bits_bridx(icache_io_cpu_btb_update_bits_prediction_bits_bridx),
    .io_cpu_btb_update_bits_prediction_bits_target(icache_io_cpu_btb_update_bits_prediction_bits_target),
    .io_cpu_btb_update_bits_prediction_bits_entry(icache_io_cpu_btb_update_bits_prediction_bits_entry),
    .io_cpu_btb_update_bits_prediction_bits_bht_history(icache_io_cpu_btb_update_bits_prediction_bits_bht_history),
    .io_cpu_btb_update_bits_prediction_bits_bht_value(icache_io_cpu_btb_update_bits_prediction_bits_bht_value),
    .io_cpu_btb_update_bits_pc(icache_io_cpu_btb_update_bits_pc),
    .io_cpu_btb_update_bits_target(icache_io_cpu_btb_update_bits_target),
    .io_cpu_btb_update_bits_taken(icache_io_cpu_btb_update_bits_taken),
    .io_cpu_btb_update_bits_isJump(icache_io_cpu_btb_update_bits_isJump),
    .io_cpu_btb_update_bits_isReturn(icache_io_cpu_btb_update_bits_isReturn),
    .io_cpu_btb_update_bits_br_pc(icache_io_cpu_btb_update_bits_br_pc),
    .io_cpu_bht_update_valid(icache_io_cpu_bht_update_valid),
    .io_cpu_bht_update_bits_prediction_valid(icache_io_cpu_bht_update_bits_prediction_valid),
    .io_cpu_bht_update_bits_prediction_bits_taken(icache_io_cpu_bht_update_bits_prediction_bits_taken),
    .io_cpu_bht_update_bits_prediction_bits_mask(icache_io_cpu_bht_update_bits_prediction_bits_mask),
    .io_cpu_bht_update_bits_prediction_bits_bridx(icache_io_cpu_bht_update_bits_prediction_bits_bridx),
    .io_cpu_bht_update_bits_prediction_bits_target(icache_io_cpu_bht_update_bits_prediction_bits_target),
    .io_cpu_bht_update_bits_prediction_bits_entry(icache_io_cpu_bht_update_bits_prediction_bits_entry),
    .io_cpu_bht_update_bits_prediction_bits_bht_history(icache_io_cpu_bht_update_bits_prediction_bits_bht_history),
    .io_cpu_bht_update_bits_prediction_bits_bht_value(icache_io_cpu_bht_update_bits_prediction_bits_bht_value),
    .io_cpu_bht_update_bits_pc(icache_io_cpu_bht_update_bits_pc),
    .io_cpu_bht_update_bits_taken(icache_io_cpu_bht_update_bits_taken),
    .io_cpu_bht_update_bits_mispredict(icache_io_cpu_bht_update_bits_mispredict),
    .io_cpu_ras_update_valid(icache_io_cpu_ras_update_valid),
    .io_cpu_ras_update_bits_isCall(icache_io_cpu_ras_update_bits_isCall),
    .io_cpu_ras_update_bits_isReturn(icache_io_cpu_ras_update_bits_isReturn),
    .io_cpu_ras_update_bits_returnAddr(icache_io_cpu_ras_update_bits_returnAddr),
    .io_cpu_ras_update_bits_prediction_valid(icache_io_cpu_ras_update_bits_prediction_valid),
    .io_cpu_ras_update_bits_prediction_bits_taken(icache_io_cpu_ras_update_bits_prediction_bits_taken),
    .io_cpu_ras_update_bits_prediction_bits_mask(icache_io_cpu_ras_update_bits_prediction_bits_mask),
    .io_cpu_ras_update_bits_prediction_bits_bridx(icache_io_cpu_ras_update_bits_prediction_bits_bridx),
    .io_cpu_ras_update_bits_prediction_bits_target(icache_io_cpu_ras_update_bits_prediction_bits_target),
    .io_cpu_ras_update_bits_prediction_bits_entry(icache_io_cpu_ras_update_bits_prediction_bits_entry),
    .io_cpu_ras_update_bits_prediction_bits_bht_history(icache_io_cpu_ras_update_bits_prediction_bits_bht_history),
    .io_cpu_ras_update_bits_prediction_bits_bht_value(icache_io_cpu_ras_update_bits_prediction_bits_bht_value),
    .io_cpu_flush_icache(icache_io_cpu_flush_icache),
    .io_cpu_flush_tlb(icache_io_cpu_flush_tlb),
    .io_cpu_npc(icache_io_cpu_npc),
    .io_ptw_req_ready(icache_io_ptw_req_ready),
    .io_ptw_req_valid(icache_io_ptw_req_valid),
    .io_ptw_req_bits_prv(icache_io_ptw_req_bits_prv),
    .io_ptw_req_bits_pum(icache_io_ptw_req_bits_pum),
    .io_ptw_req_bits_mxr(icache_io_ptw_req_bits_mxr),
    .io_ptw_req_bits_addr(icache_io_ptw_req_bits_addr),
    .io_ptw_req_bits_store(icache_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(icache_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(icache_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_reserved_for_hardware(icache_io_ptw_resp_bits_pte_reserved_for_hardware),
    .io_ptw_resp_bits_pte_ppn(icache_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(icache_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(icache_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(icache_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(icache_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(icache_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(icache_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(icache_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(icache_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(icache_io_ptw_resp_bits_pte_v),
    .io_ptw_ptbr_asid(icache_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(icache_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(icache_io_ptw_invalidate),
    .io_ptw_status_debug(icache_io_ptw_status_debug),
    .io_ptw_status_prv(icache_io_ptw_status_prv),
    .io_ptw_status_sd(icache_io_ptw_status_sd),
    .io_ptw_status_zero3(icache_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(icache_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(icache_io_ptw_status_zero2),
    .io_ptw_status_vm(icache_io_ptw_status_vm),
    .io_ptw_status_zero1(icache_io_ptw_status_zero1),
    .io_ptw_status_mxr(icache_io_ptw_status_mxr),
    .io_ptw_status_pum(icache_io_ptw_status_pum),
    .io_ptw_status_mprv(icache_io_ptw_status_mprv),
    .io_ptw_status_xs(icache_io_ptw_status_xs),
    .io_ptw_status_fs(icache_io_ptw_status_fs),
    .io_ptw_status_mpp(icache_io_ptw_status_mpp),
    .io_ptw_status_hpp(icache_io_ptw_status_hpp),
    .io_ptw_status_spp(icache_io_ptw_status_spp),
    .io_ptw_status_mpie(icache_io_ptw_status_mpie),
    .io_ptw_status_hpie(icache_io_ptw_status_hpie),
    .io_ptw_status_spie(icache_io_ptw_status_spie),
    .io_ptw_status_upie(icache_io_ptw_status_upie),
    .io_ptw_status_mie(icache_io_ptw_status_mie),
    .io_ptw_status_hie(icache_io_ptw_status_hie),
    .io_ptw_status_sie(icache_io_ptw_status_sie),
    .io_ptw_status_uie(icache_io_ptw_status_uie),
    .io_mem_acquire_ready(icache_io_mem_acquire_ready),
    .io_mem_acquire_valid(icache_io_mem_acquire_valid),
    .io_mem_acquire_bits_addr_block(icache_io_mem_acquire_bits_addr_block),
    .io_mem_acquire_bits_client_xact_id(icache_io_mem_acquire_bits_client_xact_id),
    .io_mem_acquire_bits_addr_beat(icache_io_mem_acquire_bits_addr_beat),
    .io_mem_acquire_bits_is_builtin_type(icache_io_mem_acquire_bits_is_builtin_type),
    .io_mem_acquire_bits_a_type(icache_io_mem_acquire_bits_a_type),
    .io_mem_acquire_bits_union(icache_io_mem_acquire_bits_union),
    .io_mem_acquire_bits_data(icache_io_mem_acquire_bits_data),
    .io_mem_grant_ready(icache_io_mem_grant_ready),
    .io_mem_grant_valid(icache_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(icache_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(icache_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(icache_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(icache_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(icache_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(icache_io_mem_grant_bits_data)
  );
  DCache DCache_1 (
    .clk(DCache_1_clk),
    .reset(DCache_1_reset),
    .io_cpu_req_ready(DCache_1_io_cpu_req_ready),
    .io_cpu_req_valid(DCache_1_io_cpu_req_valid),
    .io_cpu_req_bits_addr(DCache_1_io_cpu_req_bits_addr),
    .io_cpu_req_bits_tag(DCache_1_io_cpu_req_bits_tag),
    .io_cpu_req_bits_cmd(DCache_1_io_cpu_req_bits_cmd),
    .io_cpu_req_bits_typ(DCache_1_io_cpu_req_bits_typ),
    .io_cpu_req_bits_phys(DCache_1_io_cpu_req_bits_phys),
    .io_cpu_req_bits_data(DCache_1_io_cpu_req_bits_data),
    .io_cpu_s1_kill(DCache_1_io_cpu_s1_kill),
    .io_cpu_s1_data(DCache_1_io_cpu_s1_data),
    .io_cpu_s2_nack(DCache_1_io_cpu_s2_nack),
    .io_cpu_resp_valid(DCache_1_io_cpu_resp_valid),
    .io_cpu_resp_bits_addr(DCache_1_io_cpu_resp_bits_addr),
    .io_cpu_resp_bits_tag(DCache_1_io_cpu_resp_bits_tag),
    .io_cpu_resp_bits_cmd(DCache_1_io_cpu_resp_bits_cmd),
    .io_cpu_resp_bits_typ(DCache_1_io_cpu_resp_bits_typ),
    .io_cpu_resp_bits_data(DCache_1_io_cpu_resp_bits_data),
    .io_cpu_resp_bits_replay(DCache_1_io_cpu_resp_bits_replay),
    .io_cpu_resp_bits_has_data(DCache_1_io_cpu_resp_bits_has_data),
    .io_cpu_resp_bits_data_word_bypass(DCache_1_io_cpu_resp_bits_data_word_bypass),
    .io_cpu_resp_bits_store_data(DCache_1_io_cpu_resp_bits_store_data),
    .io_cpu_replay_next(DCache_1_io_cpu_replay_next),
    .io_cpu_xcpt_ma_ld(DCache_1_io_cpu_xcpt_ma_ld),
    .io_cpu_xcpt_ma_st(DCache_1_io_cpu_xcpt_ma_st),
    .io_cpu_xcpt_pf_ld(DCache_1_io_cpu_xcpt_pf_ld),
    .io_cpu_xcpt_pf_st(DCache_1_io_cpu_xcpt_pf_st),
    .io_cpu_invalidate_lr(DCache_1_io_cpu_invalidate_lr),
    .io_cpu_ordered(DCache_1_io_cpu_ordered),
    .io_ptw_req_ready(DCache_1_io_ptw_req_ready),
    .io_ptw_req_valid(DCache_1_io_ptw_req_valid),
    .io_ptw_req_bits_prv(DCache_1_io_ptw_req_bits_prv),
    .io_ptw_req_bits_pum(DCache_1_io_ptw_req_bits_pum),
    .io_ptw_req_bits_mxr(DCache_1_io_ptw_req_bits_mxr),
    .io_ptw_req_bits_addr(DCache_1_io_ptw_req_bits_addr),
    .io_ptw_req_bits_store(DCache_1_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(DCache_1_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(DCache_1_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_reserved_for_hardware(DCache_1_io_ptw_resp_bits_pte_reserved_for_hardware),
    .io_ptw_resp_bits_pte_ppn(DCache_1_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(DCache_1_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(DCache_1_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a(DCache_1_io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g(DCache_1_io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u(DCache_1_io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x(DCache_1_io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w(DCache_1_io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r(DCache_1_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v(DCache_1_io_ptw_resp_bits_pte_v),
    .io_ptw_ptbr_asid(DCache_1_io_ptw_ptbr_asid),
    .io_ptw_ptbr_ppn(DCache_1_io_ptw_ptbr_ppn),
    .io_ptw_invalidate(DCache_1_io_ptw_invalidate),
    .io_ptw_status_debug(DCache_1_io_ptw_status_debug),
    .io_ptw_status_prv(DCache_1_io_ptw_status_prv),
    .io_ptw_status_sd(DCache_1_io_ptw_status_sd),
    .io_ptw_status_zero3(DCache_1_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(DCache_1_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(DCache_1_io_ptw_status_zero2),
    .io_ptw_status_vm(DCache_1_io_ptw_status_vm),
    .io_ptw_status_zero1(DCache_1_io_ptw_status_zero1),
    .io_ptw_status_mxr(DCache_1_io_ptw_status_mxr),
    .io_ptw_status_pum(DCache_1_io_ptw_status_pum),
    .io_ptw_status_mprv(DCache_1_io_ptw_status_mprv),
    .io_ptw_status_xs(DCache_1_io_ptw_status_xs),
    .io_ptw_status_fs(DCache_1_io_ptw_status_fs),
    .io_ptw_status_mpp(DCache_1_io_ptw_status_mpp),
    .io_ptw_status_hpp(DCache_1_io_ptw_status_hpp),
    .io_ptw_status_spp(DCache_1_io_ptw_status_spp),
    .io_ptw_status_mpie(DCache_1_io_ptw_status_mpie),
    .io_ptw_status_hpie(DCache_1_io_ptw_status_hpie),
    .io_ptw_status_spie(DCache_1_io_ptw_status_spie),
    .io_ptw_status_upie(DCache_1_io_ptw_status_upie),
    .io_ptw_status_mie(DCache_1_io_ptw_status_mie),
    .io_ptw_status_hie(DCache_1_io_ptw_status_hie),
    .io_ptw_status_sie(DCache_1_io_ptw_status_sie),
    .io_ptw_status_uie(DCache_1_io_ptw_status_uie),
    .io_mem_acquire_ready(DCache_1_io_mem_acquire_ready),
    .io_mem_acquire_valid(DCache_1_io_mem_acquire_valid),
    .io_mem_acquire_bits_addr_block(DCache_1_io_mem_acquire_bits_addr_block),
    .io_mem_acquire_bits_client_xact_id(DCache_1_io_mem_acquire_bits_client_xact_id),
    .io_mem_acquire_bits_addr_beat(DCache_1_io_mem_acquire_bits_addr_beat),
    .io_mem_acquire_bits_is_builtin_type(DCache_1_io_mem_acquire_bits_is_builtin_type),
    .io_mem_acquire_bits_a_type(DCache_1_io_mem_acquire_bits_a_type),
    .io_mem_acquire_bits_union(DCache_1_io_mem_acquire_bits_union),
    .io_mem_acquire_bits_data(DCache_1_io_mem_acquire_bits_data),
    .io_mem_probe_ready(DCache_1_io_mem_probe_ready),
    .io_mem_probe_valid(DCache_1_io_mem_probe_valid),
    .io_mem_probe_bits_addr_block(DCache_1_io_mem_probe_bits_addr_block),
    .io_mem_probe_bits_p_type(DCache_1_io_mem_probe_bits_p_type),
    .io_mem_release_ready(DCache_1_io_mem_release_ready),
    .io_mem_release_valid(DCache_1_io_mem_release_valid),
    .io_mem_release_bits_addr_beat(DCache_1_io_mem_release_bits_addr_beat),
    .io_mem_release_bits_addr_block(DCache_1_io_mem_release_bits_addr_block),
    .io_mem_release_bits_client_xact_id(DCache_1_io_mem_release_bits_client_xact_id),
    .io_mem_release_bits_voluntary(DCache_1_io_mem_release_bits_voluntary),
    .io_mem_release_bits_r_type(DCache_1_io_mem_release_bits_r_type),
    .io_mem_release_bits_data(DCache_1_io_mem_release_bits_data),
    .io_mem_grant_ready(DCache_1_io_mem_grant_ready),
    .io_mem_grant_valid(DCache_1_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(DCache_1_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(DCache_1_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(DCache_1_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(DCache_1_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(DCache_1_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(DCache_1_io_mem_grant_bits_data),
    .io_mem_grant_bits_manager_id(DCache_1_io_mem_grant_bits_manager_id),
    .io_mem_finish_ready(DCache_1_io_mem_finish_ready),
    .io_mem_finish_valid(DCache_1_io_mem_finish_valid),
    .io_mem_finish_bits_manager_xact_id(DCache_1_io_mem_finish_bits_manager_xact_id),
    .io_mem_finish_bits_manager_id(DCache_1_io_mem_finish_bits_manager_id)
  );
  ClientUncachedTileLinkIOArbiter uncachedArb (
    .clk(uncachedArb_clk),
    .reset(uncachedArb_reset),
    .io_in_0_acquire_ready(uncachedArb_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(uncachedArb_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(uncachedArb_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(uncachedArb_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(uncachedArb_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(uncachedArb_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(uncachedArb_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(uncachedArb_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(uncachedArb_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(uncachedArb_io_in_0_grant_ready),
    .io_in_0_grant_valid(uncachedArb_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(uncachedArb_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(uncachedArb_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(uncachedArb_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(uncachedArb_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(uncachedArb_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(uncachedArb_io_in_0_grant_bits_data),
    .io_out_acquire_ready(uncachedArb_io_out_acquire_ready),
    .io_out_acquire_valid(uncachedArb_io_out_acquire_valid),
    .io_out_acquire_bits_addr_block(uncachedArb_io_out_acquire_bits_addr_block),
    .io_out_acquire_bits_client_xact_id(uncachedArb_io_out_acquire_bits_client_xact_id),
    .io_out_acquire_bits_addr_beat(uncachedArb_io_out_acquire_bits_addr_beat),
    .io_out_acquire_bits_is_builtin_type(uncachedArb_io_out_acquire_bits_is_builtin_type),
    .io_out_acquire_bits_a_type(uncachedArb_io_out_acquire_bits_a_type),
    .io_out_acquire_bits_union(uncachedArb_io_out_acquire_bits_union),
    .io_out_acquire_bits_data(uncachedArb_io_out_acquire_bits_data),
    .io_out_grant_ready(uncachedArb_io_out_grant_ready),
    .io_out_grant_valid(uncachedArb_io_out_grant_valid),
    .io_out_grant_bits_addr_beat(uncachedArb_io_out_grant_bits_addr_beat),
    .io_out_grant_bits_client_xact_id(uncachedArb_io_out_grant_bits_client_xact_id),
    .io_out_grant_bits_manager_xact_id(uncachedArb_io_out_grant_bits_manager_xact_id),
    .io_out_grant_bits_is_builtin_type(uncachedArb_io_out_grant_bits_is_builtin_type),
    .io_out_grant_bits_g_type(uncachedArb_io_out_grant_bits_g_type),
    .io_out_grant_bits_data(uncachedArb_io_out_grant_bits_data)
  );
  HellaCacheArbiter dcArb (
    .clk(dcArb_clk),
    .reset(dcArb_reset),
    .io_requestor_0_req_ready(dcArb_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(dcArb_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_addr(dcArb_io_requestor_0_req_bits_addr),
    .io_requestor_0_req_bits_tag(dcArb_io_requestor_0_req_bits_tag),
    .io_requestor_0_req_bits_cmd(dcArb_io_requestor_0_req_bits_cmd),
    .io_requestor_0_req_bits_typ(dcArb_io_requestor_0_req_bits_typ),
    .io_requestor_0_req_bits_phys(dcArb_io_requestor_0_req_bits_phys),
    .io_requestor_0_req_bits_data(dcArb_io_requestor_0_req_bits_data),
    .io_requestor_0_s1_kill(dcArb_io_requestor_0_s1_kill),
    .io_requestor_0_s1_data(dcArb_io_requestor_0_s1_data),
    .io_requestor_0_s2_nack(dcArb_io_requestor_0_s2_nack),
    .io_requestor_0_resp_valid(dcArb_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_addr(dcArb_io_requestor_0_resp_bits_addr),
    .io_requestor_0_resp_bits_tag(dcArb_io_requestor_0_resp_bits_tag),
    .io_requestor_0_resp_bits_cmd(dcArb_io_requestor_0_resp_bits_cmd),
    .io_requestor_0_resp_bits_typ(dcArb_io_requestor_0_resp_bits_typ),
    .io_requestor_0_resp_bits_data(dcArb_io_requestor_0_resp_bits_data),
    .io_requestor_0_resp_bits_replay(dcArb_io_requestor_0_resp_bits_replay),
    .io_requestor_0_resp_bits_has_data(dcArb_io_requestor_0_resp_bits_has_data),
    .io_requestor_0_resp_bits_data_word_bypass(dcArb_io_requestor_0_resp_bits_data_word_bypass),
    .io_requestor_0_resp_bits_store_data(dcArb_io_requestor_0_resp_bits_store_data),
    .io_requestor_0_replay_next(dcArb_io_requestor_0_replay_next),
    .io_requestor_0_xcpt_ma_ld(dcArb_io_requestor_0_xcpt_ma_ld),
    .io_requestor_0_xcpt_ma_st(dcArb_io_requestor_0_xcpt_ma_st),
    .io_requestor_0_xcpt_pf_ld(dcArb_io_requestor_0_xcpt_pf_ld),
    .io_requestor_0_xcpt_pf_st(dcArb_io_requestor_0_xcpt_pf_st),
    .io_requestor_0_invalidate_lr(dcArb_io_requestor_0_invalidate_lr),
    .io_requestor_0_ordered(dcArb_io_requestor_0_ordered),
    .io_mem_req_ready(dcArb_io_mem_req_ready),
    .io_mem_req_valid(dcArb_io_mem_req_valid),
    .io_mem_req_bits_addr(dcArb_io_mem_req_bits_addr),
    .io_mem_req_bits_tag(dcArb_io_mem_req_bits_tag),
    .io_mem_req_bits_cmd(dcArb_io_mem_req_bits_cmd),
    .io_mem_req_bits_typ(dcArb_io_mem_req_bits_typ),
    .io_mem_req_bits_phys(dcArb_io_mem_req_bits_phys),
    .io_mem_req_bits_data(dcArb_io_mem_req_bits_data),
    .io_mem_s1_kill(dcArb_io_mem_s1_kill),
    .io_mem_s1_data(dcArb_io_mem_s1_data),
    .io_mem_s2_nack(dcArb_io_mem_s2_nack),
    .io_mem_resp_valid(dcArb_io_mem_resp_valid),
    .io_mem_resp_bits_addr(dcArb_io_mem_resp_bits_addr),
    .io_mem_resp_bits_tag(dcArb_io_mem_resp_bits_tag),
    .io_mem_resp_bits_cmd(dcArb_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_typ(dcArb_io_mem_resp_bits_typ),
    .io_mem_resp_bits_data(dcArb_io_mem_resp_bits_data),
    .io_mem_resp_bits_replay(dcArb_io_mem_resp_bits_replay),
    .io_mem_resp_bits_has_data(dcArb_io_mem_resp_bits_has_data),
    .io_mem_resp_bits_data_word_bypass(dcArb_io_mem_resp_bits_data_word_bypass),
    .io_mem_resp_bits_store_data(dcArb_io_mem_resp_bits_store_data),
    .io_mem_replay_next(dcArb_io_mem_replay_next),
    .io_mem_xcpt_ma_ld(dcArb_io_mem_xcpt_ma_ld),
    .io_mem_xcpt_ma_st(dcArb_io_mem_xcpt_ma_st),
    .io_mem_xcpt_pf_ld(dcArb_io_mem_xcpt_pf_ld),
    .io_mem_xcpt_pf_st(dcArb_io_mem_xcpt_pf_st),
    .io_mem_invalidate_lr(dcArb_io_mem_invalidate_lr),
    .io_mem_ordered(dcArb_io_mem_ordered)
  );
  assign io_cached_0_acquire_valid = DCache_1_io_mem_acquire_valid;
  assign io_cached_0_acquire_bits_addr_block = DCache_1_io_mem_acquire_bits_addr_block;
  assign io_cached_0_acquire_bits_client_xact_id = DCache_1_io_mem_acquire_bits_client_xact_id;
  assign io_cached_0_acquire_bits_addr_beat = DCache_1_io_mem_acquire_bits_addr_beat;
  assign io_cached_0_acquire_bits_is_builtin_type = DCache_1_io_mem_acquire_bits_is_builtin_type;
  assign io_cached_0_acquire_bits_a_type = DCache_1_io_mem_acquire_bits_a_type;
  assign io_cached_0_acquire_bits_union = DCache_1_io_mem_acquire_bits_union;
  assign io_cached_0_acquire_bits_data = DCache_1_io_mem_acquire_bits_data;
  assign io_cached_0_probe_ready = DCache_1_io_mem_probe_ready;
  assign io_cached_0_release_valid = DCache_1_io_mem_release_valid;
  assign io_cached_0_release_bits_addr_beat = DCache_1_io_mem_release_bits_addr_beat;
  assign io_cached_0_release_bits_addr_block = DCache_1_io_mem_release_bits_addr_block;
  assign io_cached_0_release_bits_client_xact_id = DCache_1_io_mem_release_bits_client_xact_id;
  assign io_cached_0_release_bits_voluntary = DCache_1_io_mem_release_bits_voluntary;
  assign io_cached_0_release_bits_r_type = DCache_1_io_mem_release_bits_r_type;
  assign io_cached_0_release_bits_data = DCache_1_io_mem_release_bits_data;
  assign io_cached_0_grant_ready = DCache_1_io_mem_grant_ready;
  assign io_cached_0_finish_valid = DCache_1_io_mem_finish_valid;
  assign io_cached_0_finish_bits_manager_xact_id = DCache_1_io_mem_finish_bits_manager_xact_id;
  assign io_cached_0_finish_bits_manager_id = DCache_1_io_mem_finish_bits_manager_id;
  assign io_uncached_0_acquire_valid = uncachedArb_io_out_acquire_valid;
  assign io_uncached_0_acquire_bits_addr_block = uncachedArb_io_out_acquire_bits_addr_block;
  assign io_uncached_0_acquire_bits_client_xact_id = uncachedArb_io_out_acquire_bits_client_xact_id;
  assign io_uncached_0_acquire_bits_addr_beat = uncachedArb_io_out_acquire_bits_addr_beat;
  assign io_uncached_0_acquire_bits_is_builtin_type = uncachedArb_io_out_acquire_bits_is_builtin_type;
  assign io_uncached_0_acquire_bits_a_type = uncachedArb_io_out_acquire_bits_a_type;
  assign io_uncached_0_acquire_bits_union = uncachedArb_io_out_acquire_bits_union;
  assign io_uncached_0_acquire_bits_data = uncachedArb_io_out_acquire_bits_data;
  assign io_uncached_0_grant_ready = uncachedArb_io_out_grant_ready;
  assign core_clk = clk;
  assign core_reset = reset;
  assign core_io_prci_reset = io_prci_reset;
  assign core_io_prci_id = io_prci_id;
  assign core_io_prci_interrupts_meip = io_prci_interrupts_meip;
  assign core_io_prci_interrupts_seip = io_prci_interrupts_seip;
  assign core_io_prci_interrupts_debug = io_prci_interrupts_debug;
  assign core_io_prci_interrupts_mtip = io_prci_interrupts_mtip;
  assign core_io_prci_interrupts_msip = io_prci_interrupts_msip;
  assign core_io_imem_resp_valid = icache_io_cpu_resp_valid;
  assign core_io_imem_resp_bits_pc = icache_io_cpu_resp_bits_pc;
  assign core_io_imem_resp_bits_data_0 = icache_io_cpu_resp_bits_data_0;
  assign core_io_imem_resp_bits_mask = icache_io_cpu_resp_bits_mask;
  assign core_io_imem_resp_bits_xcpt_if = icache_io_cpu_resp_bits_xcpt_if;
  assign core_io_imem_resp_bits_replay = icache_io_cpu_resp_bits_replay;
  assign core_io_imem_btb_resp_valid = icache_io_cpu_btb_resp_valid;
  assign core_io_imem_btb_resp_bits_taken = icache_io_cpu_btb_resp_bits_taken;
  assign core_io_imem_btb_resp_bits_mask = icache_io_cpu_btb_resp_bits_mask;
  assign core_io_imem_btb_resp_bits_bridx = icache_io_cpu_btb_resp_bits_bridx;
  assign core_io_imem_btb_resp_bits_target = icache_io_cpu_btb_resp_bits_target;
  assign core_io_imem_btb_resp_bits_entry = icache_io_cpu_btb_resp_bits_entry;
  assign core_io_imem_btb_resp_bits_bht_history = icache_io_cpu_btb_resp_bits_bht_history;
  assign core_io_imem_btb_resp_bits_bht_value = icache_io_cpu_btb_resp_bits_bht_value;
  assign core_io_imem_npc = icache_io_cpu_npc;
  assign core_io_dmem_req_ready = dcArb_io_requestor_0_req_ready;
  assign core_io_dmem_s2_nack = dcArb_io_requestor_0_s2_nack;
  assign core_io_dmem_resp_valid = dcArb_io_requestor_0_resp_valid;
  assign core_io_dmem_resp_bits_addr = dcArb_io_requestor_0_resp_bits_addr;
  assign core_io_dmem_resp_bits_tag = dcArb_io_requestor_0_resp_bits_tag;
  assign core_io_dmem_resp_bits_cmd = dcArb_io_requestor_0_resp_bits_cmd;
  assign core_io_dmem_resp_bits_typ = dcArb_io_requestor_0_resp_bits_typ;
  assign core_io_dmem_resp_bits_data = dcArb_io_requestor_0_resp_bits_data;
  assign core_io_dmem_resp_bits_replay = dcArb_io_requestor_0_resp_bits_replay;
  assign core_io_dmem_resp_bits_has_data = dcArb_io_requestor_0_resp_bits_has_data;
  assign core_io_dmem_resp_bits_data_word_bypass = dcArb_io_requestor_0_resp_bits_data_word_bypass;
  assign core_io_dmem_resp_bits_store_data = dcArb_io_requestor_0_resp_bits_store_data;
  assign core_io_dmem_replay_next = dcArb_io_requestor_0_replay_next;
  assign core_io_dmem_xcpt_ma_ld = dcArb_io_requestor_0_xcpt_ma_ld;
  assign core_io_dmem_xcpt_ma_st = dcArb_io_requestor_0_xcpt_ma_st;
  assign core_io_dmem_xcpt_pf_ld = dcArb_io_requestor_0_xcpt_pf_ld;
  assign core_io_dmem_xcpt_pf_st = dcArb_io_requestor_0_xcpt_pf_st;
  assign core_io_dmem_ordered = dcArb_io_requestor_0_ordered;
  assign core_io_fpu_fcsr_flags_valid = GEN_0;
  assign core_io_fpu_fcsr_flags_bits = GEN_1;
  assign core_io_fpu_store_data = GEN_2;
  assign core_io_fpu_toint_data = GEN_3;
  assign core_io_fpu_fcsr_rdy = GEN_4;
  assign core_io_fpu_nack_mem = GEN_5;
  assign core_io_fpu_illegal_rm = GEN_6;
  assign core_io_fpu_dec_cmd = GEN_7;
  assign core_io_fpu_dec_ldst = GEN_8;
  assign core_io_fpu_dec_wen = GEN_9;
  assign core_io_fpu_dec_ren1 = GEN_10;
  assign core_io_fpu_dec_ren2 = GEN_11;
  assign core_io_fpu_dec_ren3 = GEN_12;
  assign core_io_fpu_dec_swap12 = GEN_13;
  assign core_io_fpu_dec_swap23 = GEN_14;
  assign core_io_fpu_dec_single = GEN_15;
  assign core_io_fpu_dec_fromint = GEN_16;
  assign core_io_fpu_dec_toint = GEN_17;
  assign core_io_fpu_dec_fastpipe = GEN_18;
  assign core_io_fpu_dec_fma = GEN_19;
  assign core_io_fpu_dec_div = GEN_20;
  assign core_io_fpu_dec_sqrt = GEN_21;
  assign core_io_fpu_dec_round = GEN_22;
  assign core_io_fpu_dec_wflags = GEN_23;
  assign core_io_fpu_sboard_set = GEN_24;
  assign core_io_fpu_sboard_clr = GEN_25;
  assign core_io_fpu_sboard_clra = GEN_26;
  assign core_io_fpu_cp_req_ready = GEN_27;
  assign core_io_fpu_cp_resp_valid = GEN_28;
  assign core_io_fpu_cp_resp_bits_data = GEN_29;
  assign core_io_fpu_cp_resp_bits_exc = GEN_30;
  assign core_io_rocc_cmd_ready = GEN_31;
  assign core_io_rocc_resp_valid = GEN_32;
  assign core_io_rocc_resp_bits_rd = GEN_33;
  assign core_io_rocc_resp_bits_data = GEN_34;
  assign core_io_rocc_mem_req_valid = GEN_35;
  assign core_io_rocc_mem_req_bits_addr = GEN_36;
  assign core_io_rocc_mem_req_bits_tag = GEN_37;
  assign core_io_rocc_mem_req_bits_cmd = GEN_38;
  assign core_io_rocc_mem_req_bits_typ = GEN_39;
  assign core_io_rocc_mem_req_bits_phys = GEN_40;
  assign core_io_rocc_mem_req_bits_data = GEN_41;
  assign core_io_rocc_mem_s1_kill = GEN_42;
  assign core_io_rocc_mem_s1_data = GEN_43;
  assign core_io_rocc_mem_invalidate_lr = GEN_44;
  assign core_io_rocc_busy = GEN_45;
  assign core_io_rocc_interrupt = GEN_46;
  assign core_io_rocc_autl_acquire_valid = GEN_47;
  assign core_io_rocc_autl_acquire_bits_addr_block = GEN_48;
  assign core_io_rocc_autl_acquire_bits_client_xact_id = GEN_49;
  assign core_io_rocc_autl_acquire_bits_addr_beat = GEN_50;
  assign core_io_rocc_autl_acquire_bits_is_builtin_type = GEN_51;
  assign core_io_rocc_autl_acquire_bits_a_type = GEN_52;
  assign core_io_rocc_autl_acquire_bits_union = GEN_53;
  assign core_io_rocc_autl_acquire_bits_data = GEN_54;
  assign core_io_rocc_autl_grant_ready = GEN_55;
  assign core_io_rocc_fpu_req_valid = GEN_56;
  assign core_io_rocc_fpu_req_bits_cmd = GEN_57;
  assign core_io_rocc_fpu_req_bits_ldst = GEN_58;
  assign core_io_rocc_fpu_req_bits_wen = GEN_59;
  assign core_io_rocc_fpu_req_bits_ren1 = GEN_60;
  assign core_io_rocc_fpu_req_bits_ren2 = GEN_61;
  assign core_io_rocc_fpu_req_bits_ren3 = GEN_62;
  assign core_io_rocc_fpu_req_bits_swap12 = GEN_63;
  assign core_io_rocc_fpu_req_bits_swap23 = GEN_64;
  assign core_io_rocc_fpu_req_bits_single = GEN_65;
  assign core_io_rocc_fpu_req_bits_fromint = GEN_66;
  assign core_io_rocc_fpu_req_bits_toint = GEN_67;
  assign core_io_rocc_fpu_req_bits_fastpipe = GEN_68;
  assign core_io_rocc_fpu_req_bits_fma = GEN_69;
  assign core_io_rocc_fpu_req_bits_div = GEN_70;
  assign core_io_rocc_fpu_req_bits_sqrt = GEN_71;
  assign core_io_rocc_fpu_req_bits_round = GEN_72;
  assign core_io_rocc_fpu_req_bits_wflags = GEN_73;
  assign core_io_rocc_fpu_req_bits_rm = GEN_74;
  assign core_io_rocc_fpu_req_bits_typ = GEN_75;
  assign core_io_rocc_fpu_req_bits_in1 = GEN_76;
  assign core_io_rocc_fpu_req_bits_in2 = GEN_77;
  assign core_io_rocc_fpu_req_bits_in3 = GEN_78;
  assign core_io_rocc_fpu_resp_ready = GEN_79;
  assign icache_clk = clk;
  assign icache_reset = reset;
  assign icache_io_cpu_req_valid = core_io_imem_req_valid;
  assign icache_io_cpu_req_bits_pc = core_io_imem_req_bits_pc;
  assign icache_io_cpu_req_bits_speculative = core_io_imem_req_bits_speculative;
  assign icache_io_cpu_resp_ready = core_io_imem_resp_ready;
  assign icache_io_cpu_btb_update_valid = core_io_imem_btb_update_valid;
  assign icache_io_cpu_btb_update_bits_prediction_valid = core_io_imem_btb_update_bits_prediction_valid;
  assign icache_io_cpu_btb_update_bits_prediction_bits_taken = core_io_imem_btb_update_bits_prediction_bits_taken;
  assign icache_io_cpu_btb_update_bits_prediction_bits_mask = core_io_imem_btb_update_bits_prediction_bits_mask;
  assign icache_io_cpu_btb_update_bits_prediction_bits_bridx = core_io_imem_btb_update_bits_prediction_bits_bridx;
  assign icache_io_cpu_btb_update_bits_prediction_bits_target = core_io_imem_btb_update_bits_prediction_bits_target;
  assign icache_io_cpu_btb_update_bits_prediction_bits_entry = core_io_imem_btb_update_bits_prediction_bits_entry;
  assign icache_io_cpu_btb_update_bits_prediction_bits_bht_history = core_io_imem_btb_update_bits_prediction_bits_bht_history;
  assign icache_io_cpu_btb_update_bits_prediction_bits_bht_value = core_io_imem_btb_update_bits_prediction_bits_bht_value;
  assign icache_io_cpu_btb_update_bits_pc = core_io_imem_btb_update_bits_pc;
  assign icache_io_cpu_btb_update_bits_target = core_io_imem_btb_update_bits_target;
  assign icache_io_cpu_btb_update_bits_taken = core_io_imem_btb_update_bits_taken;
  assign icache_io_cpu_btb_update_bits_isJump = core_io_imem_btb_update_bits_isJump;
  assign icache_io_cpu_btb_update_bits_isReturn = core_io_imem_btb_update_bits_isReturn;
  assign icache_io_cpu_btb_update_bits_br_pc = core_io_imem_btb_update_bits_br_pc;
  assign icache_io_cpu_bht_update_valid = core_io_imem_bht_update_valid;
  assign icache_io_cpu_bht_update_bits_prediction_valid = core_io_imem_bht_update_bits_prediction_valid;
  assign icache_io_cpu_bht_update_bits_prediction_bits_taken = core_io_imem_bht_update_bits_prediction_bits_taken;
  assign icache_io_cpu_bht_update_bits_prediction_bits_mask = core_io_imem_bht_update_bits_prediction_bits_mask;
  assign icache_io_cpu_bht_update_bits_prediction_bits_bridx = core_io_imem_bht_update_bits_prediction_bits_bridx;
  assign icache_io_cpu_bht_update_bits_prediction_bits_target = core_io_imem_bht_update_bits_prediction_bits_target;
  assign icache_io_cpu_bht_update_bits_prediction_bits_entry = core_io_imem_bht_update_bits_prediction_bits_entry;
  assign icache_io_cpu_bht_update_bits_prediction_bits_bht_history = core_io_imem_bht_update_bits_prediction_bits_bht_history;
  assign icache_io_cpu_bht_update_bits_prediction_bits_bht_value = core_io_imem_bht_update_bits_prediction_bits_bht_value;
  assign icache_io_cpu_bht_update_bits_pc = core_io_imem_bht_update_bits_pc;
  assign icache_io_cpu_bht_update_bits_taken = core_io_imem_bht_update_bits_taken;
  assign icache_io_cpu_bht_update_bits_mispredict = core_io_imem_bht_update_bits_mispredict;
  assign icache_io_cpu_ras_update_valid = core_io_imem_ras_update_valid;
  assign icache_io_cpu_ras_update_bits_isCall = core_io_imem_ras_update_bits_isCall;
  assign icache_io_cpu_ras_update_bits_isReturn = core_io_imem_ras_update_bits_isReturn;
  assign icache_io_cpu_ras_update_bits_returnAddr = core_io_imem_ras_update_bits_returnAddr;
  assign icache_io_cpu_ras_update_bits_prediction_valid = core_io_imem_ras_update_bits_prediction_valid;
  assign icache_io_cpu_ras_update_bits_prediction_bits_taken = core_io_imem_ras_update_bits_prediction_bits_taken;
  assign icache_io_cpu_ras_update_bits_prediction_bits_mask = core_io_imem_ras_update_bits_prediction_bits_mask;
  assign icache_io_cpu_ras_update_bits_prediction_bits_bridx = core_io_imem_ras_update_bits_prediction_bits_bridx;
  assign icache_io_cpu_ras_update_bits_prediction_bits_target = core_io_imem_ras_update_bits_prediction_bits_target;
  assign icache_io_cpu_ras_update_bits_prediction_bits_entry = core_io_imem_ras_update_bits_prediction_bits_entry;
  assign icache_io_cpu_ras_update_bits_prediction_bits_bht_history = core_io_imem_ras_update_bits_prediction_bits_bht_history;
  assign icache_io_cpu_ras_update_bits_prediction_bits_bht_value = core_io_imem_ras_update_bits_prediction_bits_bht_value;
  assign icache_io_cpu_flush_icache = core_io_imem_flush_icache;
  assign icache_io_cpu_flush_tlb = core_io_imem_flush_tlb;
  assign icache_io_ptw_req_ready = GEN_80;
  assign icache_io_ptw_resp_valid = GEN_81;
  assign icache_io_ptw_resp_bits_pte_reserved_for_hardware = GEN_82;
  assign icache_io_ptw_resp_bits_pte_ppn = GEN_83;
  assign icache_io_ptw_resp_bits_pte_reserved_for_software = GEN_84;
  assign icache_io_ptw_resp_bits_pte_d = GEN_85;
  assign icache_io_ptw_resp_bits_pte_a = GEN_86;
  assign icache_io_ptw_resp_bits_pte_g = GEN_87;
  assign icache_io_ptw_resp_bits_pte_u = GEN_88;
  assign icache_io_ptw_resp_bits_pte_x = GEN_89;
  assign icache_io_ptw_resp_bits_pte_w = GEN_90;
  assign icache_io_ptw_resp_bits_pte_r = GEN_91;
  assign icache_io_ptw_resp_bits_pte_v = GEN_92;
  assign icache_io_ptw_ptbr_asid = GEN_93;
  assign icache_io_ptw_ptbr_ppn = GEN_94;
  assign icache_io_ptw_invalidate = GEN_95;
  assign icache_io_ptw_status_debug = GEN_96;
  assign icache_io_ptw_status_prv = GEN_97;
  assign icache_io_ptw_status_sd = GEN_98;
  assign icache_io_ptw_status_zero3 = GEN_99;
  assign icache_io_ptw_status_sd_rv32 = GEN_100;
  assign icache_io_ptw_status_zero2 = GEN_101;
  assign icache_io_ptw_status_vm = GEN_102;
  assign icache_io_ptw_status_zero1 = GEN_103;
  assign icache_io_ptw_status_mxr = GEN_104;
  assign icache_io_ptw_status_pum = GEN_105;
  assign icache_io_ptw_status_mprv = GEN_106;
  assign icache_io_ptw_status_xs = GEN_107;
  assign icache_io_ptw_status_fs = GEN_108;
  assign icache_io_ptw_status_mpp = GEN_109;
  assign icache_io_ptw_status_hpp = GEN_110;
  assign icache_io_ptw_status_spp = GEN_111;
  assign icache_io_ptw_status_mpie = GEN_112;
  assign icache_io_ptw_status_hpie = GEN_113;
  assign icache_io_ptw_status_spie = GEN_114;
  assign icache_io_ptw_status_upie = GEN_115;
  assign icache_io_ptw_status_mie = GEN_116;
  assign icache_io_ptw_status_hie = GEN_117;
  assign icache_io_ptw_status_sie = GEN_118;
  assign icache_io_ptw_status_uie = GEN_119;
  assign icache_io_mem_acquire_ready = uncachedArb_io_in_0_acquire_ready;
  assign icache_io_mem_grant_valid = uncachedArb_io_in_0_grant_valid;
  assign icache_io_mem_grant_bits_addr_beat = uncachedArb_io_in_0_grant_bits_addr_beat;
  assign icache_io_mem_grant_bits_client_xact_id = uncachedArb_io_in_0_grant_bits_client_xact_id;
  assign icache_io_mem_grant_bits_manager_xact_id = uncachedArb_io_in_0_grant_bits_manager_xact_id;
  assign icache_io_mem_grant_bits_is_builtin_type = uncachedArb_io_in_0_grant_bits_is_builtin_type;
  assign icache_io_mem_grant_bits_g_type = uncachedArb_io_in_0_grant_bits_g_type;
  assign icache_io_mem_grant_bits_data = uncachedArb_io_in_0_grant_bits_data;
  assign DCache_1_clk = clk;
  assign DCache_1_reset = reset;
  assign DCache_1_io_cpu_req_valid = dcArb_io_mem_req_valid;
  assign DCache_1_io_cpu_req_bits_addr = dcArb_io_mem_req_bits_addr;
  assign DCache_1_io_cpu_req_bits_tag = dcArb_io_mem_req_bits_tag;
  assign DCache_1_io_cpu_req_bits_cmd = dcArb_io_mem_req_bits_cmd;
  assign DCache_1_io_cpu_req_bits_typ = dcArb_io_mem_req_bits_typ;
  assign DCache_1_io_cpu_req_bits_phys = dcArb_io_mem_req_bits_phys;
  assign DCache_1_io_cpu_req_bits_data = dcArb_io_mem_req_bits_data;
  assign DCache_1_io_cpu_s1_kill = dcArb_io_mem_s1_kill;
  assign DCache_1_io_cpu_s1_data = dcArb_io_mem_s1_data;
  assign DCache_1_io_cpu_invalidate_lr = dcArb_io_mem_invalidate_lr;
  assign DCache_1_io_ptw_req_ready = GEN_120;
  assign DCache_1_io_ptw_resp_valid = GEN_121;
  assign DCache_1_io_ptw_resp_bits_pte_reserved_for_hardware = GEN_122;
  assign DCache_1_io_ptw_resp_bits_pte_ppn = GEN_123;
  assign DCache_1_io_ptw_resp_bits_pte_reserved_for_software = GEN_124;
  assign DCache_1_io_ptw_resp_bits_pte_d = GEN_125;
  assign DCache_1_io_ptw_resp_bits_pte_a = GEN_126;
  assign DCache_1_io_ptw_resp_bits_pte_g = GEN_127;
  assign DCache_1_io_ptw_resp_bits_pte_u = GEN_128;
  assign DCache_1_io_ptw_resp_bits_pte_x = GEN_129;
  assign DCache_1_io_ptw_resp_bits_pte_w = GEN_130;
  assign DCache_1_io_ptw_resp_bits_pte_r = GEN_131;
  assign DCache_1_io_ptw_resp_bits_pte_v = GEN_132;
  assign DCache_1_io_ptw_ptbr_asid = GEN_133;
  assign DCache_1_io_ptw_ptbr_ppn = GEN_134;
  assign DCache_1_io_ptw_invalidate = GEN_135;
  assign DCache_1_io_ptw_status_debug = GEN_136;
  assign DCache_1_io_ptw_status_prv = GEN_137;
  assign DCache_1_io_ptw_status_sd = GEN_138;
  assign DCache_1_io_ptw_status_zero3 = GEN_139;
  assign DCache_1_io_ptw_status_sd_rv32 = GEN_140;
  assign DCache_1_io_ptw_status_zero2 = GEN_141;
  assign DCache_1_io_ptw_status_vm = GEN_142;
  assign DCache_1_io_ptw_status_zero1 = GEN_143;
  assign DCache_1_io_ptw_status_mxr = GEN_144;
  assign DCache_1_io_ptw_status_pum = GEN_145;
  assign DCache_1_io_ptw_status_mprv = GEN_146;
  assign DCache_1_io_ptw_status_xs = GEN_147;
  assign DCache_1_io_ptw_status_fs = GEN_148;
  assign DCache_1_io_ptw_status_mpp = GEN_149;
  assign DCache_1_io_ptw_status_hpp = GEN_150;
  assign DCache_1_io_ptw_status_spp = GEN_151;
  assign DCache_1_io_ptw_status_mpie = GEN_152;
  assign DCache_1_io_ptw_status_hpie = GEN_153;
  assign DCache_1_io_ptw_status_spie = GEN_154;
  assign DCache_1_io_ptw_status_upie = GEN_155;
  assign DCache_1_io_ptw_status_mie = GEN_156;
  assign DCache_1_io_ptw_status_hie = GEN_157;
  assign DCache_1_io_ptw_status_sie = GEN_158;
  assign DCache_1_io_ptw_status_uie = GEN_159;
  assign DCache_1_io_mem_acquire_ready = io_cached_0_acquire_ready;
  assign DCache_1_io_mem_probe_valid = io_cached_0_probe_valid;
  assign DCache_1_io_mem_probe_bits_addr_block = io_cached_0_probe_bits_addr_block;
  assign DCache_1_io_mem_probe_bits_p_type = io_cached_0_probe_bits_p_type;
  assign DCache_1_io_mem_release_ready = io_cached_0_release_ready;
  assign DCache_1_io_mem_grant_valid = io_cached_0_grant_valid;
  assign DCache_1_io_mem_grant_bits_addr_beat = io_cached_0_grant_bits_addr_beat;
  assign DCache_1_io_mem_grant_bits_client_xact_id = io_cached_0_grant_bits_client_xact_id;
  assign DCache_1_io_mem_grant_bits_manager_xact_id = io_cached_0_grant_bits_manager_xact_id;
  assign DCache_1_io_mem_grant_bits_is_builtin_type = io_cached_0_grant_bits_is_builtin_type;
  assign DCache_1_io_mem_grant_bits_g_type = io_cached_0_grant_bits_g_type;
  assign DCache_1_io_mem_grant_bits_data = io_cached_0_grant_bits_data;
  assign DCache_1_io_mem_grant_bits_manager_id = io_cached_0_grant_bits_manager_id;
  assign DCache_1_io_mem_finish_ready = io_cached_0_finish_ready;
  assign uncachedArb_clk = clk;
  assign uncachedArb_reset = reset;
  assign uncachedArb_io_in_0_acquire_valid = icache_io_mem_acquire_valid;
  assign uncachedArb_io_in_0_acquire_bits_addr_block = icache_io_mem_acquire_bits_addr_block;
  assign uncachedArb_io_in_0_acquire_bits_client_xact_id = icache_io_mem_acquire_bits_client_xact_id;
  assign uncachedArb_io_in_0_acquire_bits_addr_beat = icache_io_mem_acquire_bits_addr_beat;
  assign uncachedArb_io_in_0_acquire_bits_is_builtin_type = icache_io_mem_acquire_bits_is_builtin_type;
  assign uncachedArb_io_in_0_acquire_bits_a_type = icache_io_mem_acquire_bits_a_type;
  assign uncachedArb_io_in_0_acquire_bits_union = icache_io_mem_acquire_bits_union;
  assign uncachedArb_io_in_0_acquire_bits_data = icache_io_mem_acquire_bits_data;
  assign uncachedArb_io_in_0_grant_ready = icache_io_mem_grant_ready;
  assign uncachedArb_io_out_acquire_ready = io_uncached_0_acquire_ready;
  assign uncachedArb_io_out_grant_valid = io_uncached_0_grant_valid;
  assign uncachedArb_io_out_grant_bits_addr_beat = io_uncached_0_grant_bits_addr_beat;
  assign uncachedArb_io_out_grant_bits_client_xact_id = io_uncached_0_grant_bits_client_xact_id;
  assign uncachedArb_io_out_grant_bits_manager_xact_id = io_uncached_0_grant_bits_manager_xact_id;
  assign uncachedArb_io_out_grant_bits_is_builtin_type = io_uncached_0_grant_bits_is_builtin_type;
  assign uncachedArb_io_out_grant_bits_g_type = io_uncached_0_grant_bits_g_type;
  assign uncachedArb_io_out_grant_bits_data = io_uncached_0_grant_bits_data;
  assign dcArb_clk = clk;
  assign dcArb_reset = reset;
  assign dcArb_io_requestor_0_req_valid = core_io_dmem_req_valid;
  assign dcArb_io_requestor_0_req_bits_addr = core_io_dmem_req_bits_addr;
  assign dcArb_io_requestor_0_req_bits_tag = core_io_dmem_req_bits_tag;
  assign dcArb_io_requestor_0_req_bits_cmd = core_io_dmem_req_bits_cmd;
  assign dcArb_io_requestor_0_req_bits_typ = core_io_dmem_req_bits_typ;
  assign dcArb_io_requestor_0_req_bits_phys = core_io_dmem_req_bits_phys;
  assign dcArb_io_requestor_0_req_bits_data = core_io_dmem_req_bits_data;
  assign dcArb_io_requestor_0_s1_kill = core_io_dmem_s1_kill;
  assign dcArb_io_requestor_0_s1_data = core_io_dmem_s1_data;
  assign dcArb_io_requestor_0_invalidate_lr = core_io_dmem_invalidate_lr;
  assign dcArb_io_mem_req_ready = DCache_1_io_cpu_req_ready;
  assign dcArb_io_mem_s2_nack = DCache_1_io_cpu_s2_nack;
  assign dcArb_io_mem_resp_valid = DCache_1_io_cpu_resp_valid;
  assign dcArb_io_mem_resp_bits_addr = DCache_1_io_cpu_resp_bits_addr;
  assign dcArb_io_mem_resp_bits_tag = DCache_1_io_cpu_resp_bits_tag;
  assign dcArb_io_mem_resp_bits_cmd = DCache_1_io_cpu_resp_bits_cmd;
  assign dcArb_io_mem_resp_bits_typ = DCache_1_io_cpu_resp_bits_typ;
  assign dcArb_io_mem_resp_bits_data = DCache_1_io_cpu_resp_bits_data;
  assign dcArb_io_mem_resp_bits_replay = DCache_1_io_cpu_resp_bits_replay;
  assign dcArb_io_mem_resp_bits_has_data = DCache_1_io_cpu_resp_bits_has_data;
  assign dcArb_io_mem_resp_bits_data_word_bypass = DCache_1_io_cpu_resp_bits_data_word_bypass;
  assign dcArb_io_mem_resp_bits_store_data = DCache_1_io_cpu_resp_bits_store_data;
  assign dcArb_io_mem_replay_next = DCache_1_io_cpu_replay_next;
  assign dcArb_io_mem_xcpt_ma_ld = DCache_1_io_cpu_xcpt_ma_ld;
  assign dcArb_io_mem_xcpt_ma_st = DCache_1_io_cpu_xcpt_ma_st;
  assign dcArb_io_mem_xcpt_pf_ld = DCache_1_io_cpu_xcpt_pf_ld;
  assign dcArb_io_mem_xcpt_pf_st = DCache_1_io_cpu_xcpt_pf_st;
  assign dcArb_io_mem_ordered = DCache_1_io_cpu_ordered;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_160 = {1{$random}};
  GEN_0 = GEN_160[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_161 = {1{$random}};
  GEN_1 = GEN_161[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_162 = {2{$random}};
  GEN_2 = GEN_162[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_163 = {1{$random}};
  GEN_3 = GEN_163[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_164 = {1{$random}};
  GEN_4 = GEN_164[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_165 = {1{$random}};
  GEN_5 = GEN_165[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_166 = {1{$random}};
  GEN_6 = GEN_166[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_167 = {1{$random}};
  GEN_7 = GEN_167[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_168 = {1{$random}};
  GEN_8 = GEN_168[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_169 = {1{$random}};
  GEN_9 = GEN_169[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_170 = {1{$random}};
  GEN_10 = GEN_170[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_171 = {1{$random}};
  GEN_11 = GEN_171[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_172 = {1{$random}};
  GEN_12 = GEN_172[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_173 = {1{$random}};
  GEN_13 = GEN_173[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_174 = {1{$random}};
  GEN_14 = GEN_174[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_175 = {1{$random}};
  GEN_15 = GEN_175[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_176 = {1{$random}};
  GEN_16 = GEN_176[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_177 = {1{$random}};
  GEN_17 = GEN_177[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_178 = {1{$random}};
  GEN_18 = GEN_178[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_179 = {1{$random}};
  GEN_19 = GEN_179[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_180 = {1{$random}};
  GEN_20 = GEN_180[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_181 = {1{$random}};
  GEN_21 = GEN_181[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_182 = {1{$random}};
  GEN_22 = GEN_182[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_183 = {1{$random}};
  GEN_23 = GEN_183[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_184 = {1{$random}};
  GEN_24 = GEN_184[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_185 = {1{$random}};
  GEN_25 = GEN_185[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_186 = {1{$random}};
  GEN_26 = GEN_186[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_187 = {1{$random}};
  GEN_27 = GEN_187[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_188 = {1{$random}};
  GEN_28 = GEN_188[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_189 = {3{$random}};
  GEN_29 = GEN_189[64:0];
  `endif
  `ifdef RANDOMIZE
  GEN_190 = {1{$random}};
  GEN_30 = GEN_190[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_191 = {1{$random}};
  GEN_31 = GEN_191[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_192 = {1{$random}};
  GEN_32 = GEN_192[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_193 = {1{$random}};
  GEN_33 = GEN_193[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_194 = {1{$random}};
  GEN_34 = GEN_194[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_195 = {1{$random}};
  GEN_35 = GEN_195[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_196 = {1{$random}};
  GEN_36 = GEN_196[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_197 = {1{$random}};
  GEN_37 = GEN_197[8:0];
  `endif
  `ifdef RANDOMIZE
  GEN_198 = {1{$random}};
  GEN_38 = GEN_198[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_199 = {1{$random}};
  GEN_39 = GEN_199[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_200 = {1{$random}};
  GEN_40 = GEN_200[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_201 = {1{$random}};
  GEN_41 = GEN_201[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_202 = {1{$random}};
  GEN_42 = GEN_202[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_203 = {1{$random}};
  GEN_43 = GEN_203[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_204 = {1{$random}};
  GEN_44 = GEN_204[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_205 = {1{$random}};
  GEN_45 = GEN_205[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_206 = {1{$random}};
  GEN_46 = GEN_206[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_207 = {1{$random}};
  GEN_47 = GEN_207[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_208 = {1{$random}};
  GEN_48 = GEN_208[25:0];
  `endif
  `ifdef RANDOMIZE
  GEN_209 = {1{$random}};
  GEN_49 = GEN_209[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_210 = {1{$random}};
  GEN_50 = GEN_210[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_211 = {1{$random}};
  GEN_51 = GEN_211[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_212 = {1{$random}};
  GEN_52 = GEN_212[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_213 = {1{$random}};
  GEN_53 = GEN_213[11:0];
  `endif
  `ifdef RANDOMIZE
  GEN_214 = {2{$random}};
  GEN_54 = GEN_214[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_215 = {1{$random}};
  GEN_55 = GEN_215[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_216 = {1{$random}};
  GEN_56 = GEN_216[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_217 = {1{$random}};
  GEN_57 = GEN_217[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_218 = {1{$random}};
  GEN_58 = GEN_218[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_219 = {1{$random}};
  GEN_59 = GEN_219[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_220 = {1{$random}};
  GEN_60 = GEN_220[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_221 = {1{$random}};
  GEN_61 = GEN_221[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_222 = {1{$random}};
  GEN_62 = GEN_222[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_223 = {1{$random}};
  GEN_63 = GEN_223[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_224 = {1{$random}};
  GEN_64 = GEN_224[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_225 = {1{$random}};
  GEN_65 = GEN_225[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_226 = {1{$random}};
  GEN_66 = GEN_226[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_227 = {1{$random}};
  GEN_67 = GEN_227[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_228 = {1{$random}};
  GEN_68 = GEN_228[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_229 = {1{$random}};
  GEN_69 = GEN_229[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_230 = {1{$random}};
  GEN_70 = GEN_230[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_231 = {1{$random}};
  GEN_71 = GEN_231[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_232 = {1{$random}};
  GEN_72 = GEN_232[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_233 = {1{$random}};
  GEN_73 = GEN_233[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_234 = {1{$random}};
  GEN_74 = GEN_234[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_235 = {1{$random}};
  GEN_75 = GEN_235[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_236 = {3{$random}};
  GEN_76 = GEN_236[64:0];
  `endif
  `ifdef RANDOMIZE
  GEN_237 = {3{$random}};
  GEN_77 = GEN_237[64:0];
  `endif
  `ifdef RANDOMIZE
  GEN_238 = {3{$random}};
  GEN_78 = GEN_238[64:0];
  `endif
  `ifdef RANDOMIZE
  GEN_239 = {1{$random}};
  GEN_79 = GEN_239[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_240 = {1{$random}};
  GEN_80 = GEN_240[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_241 = {1{$random}};
  GEN_81 = GEN_241[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_242 = {1{$random}};
  GEN_82 = GEN_242[15:0];
  `endif
  `ifdef RANDOMIZE
  GEN_243 = {2{$random}};
  GEN_83 = GEN_243[37:0];
  `endif
  `ifdef RANDOMIZE
  GEN_244 = {1{$random}};
  GEN_84 = GEN_244[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_245 = {1{$random}};
  GEN_85 = GEN_245[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_246 = {1{$random}};
  GEN_86 = GEN_246[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_247 = {1{$random}};
  GEN_87 = GEN_247[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_248 = {1{$random}};
  GEN_88 = GEN_248[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_249 = {1{$random}};
  GEN_89 = GEN_249[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_250 = {1{$random}};
  GEN_90 = GEN_250[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_251 = {1{$random}};
  GEN_91 = GEN_251[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_252 = {1{$random}};
  GEN_92 = GEN_252[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_253 = {1{$random}};
  GEN_93 = GEN_253[6:0];
  `endif
  `ifdef RANDOMIZE
  GEN_254 = {1{$random}};
  GEN_94 = GEN_254[21:0];
  `endif
  `ifdef RANDOMIZE
  GEN_255 = {1{$random}};
  GEN_95 = GEN_255[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_256 = {1{$random}};
  GEN_96 = GEN_256[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_257 = {1{$random}};
  GEN_97 = GEN_257[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_258 = {1{$random}};
  GEN_98 = GEN_258[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_259 = {1{$random}};
  GEN_99 = GEN_259[30:0];
  `endif
  `ifdef RANDOMIZE
  GEN_260 = {1{$random}};
  GEN_100 = GEN_260[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_261 = {1{$random}};
  GEN_101 = GEN_261[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_262 = {1{$random}};
  GEN_102 = GEN_262[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_263 = {1{$random}};
  GEN_103 = GEN_263[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_264 = {1{$random}};
  GEN_104 = GEN_264[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_265 = {1{$random}};
  GEN_105 = GEN_265[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_266 = {1{$random}};
  GEN_106 = GEN_266[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_267 = {1{$random}};
  GEN_107 = GEN_267[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_268 = {1{$random}};
  GEN_108 = GEN_268[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_269 = {1{$random}};
  GEN_109 = GEN_269[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_270 = {1{$random}};
  GEN_110 = GEN_270[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_271 = {1{$random}};
  GEN_111 = GEN_271[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_272 = {1{$random}};
  GEN_112 = GEN_272[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_273 = {1{$random}};
  GEN_113 = GEN_273[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_274 = {1{$random}};
  GEN_114 = GEN_274[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_275 = {1{$random}};
  GEN_115 = GEN_275[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_276 = {1{$random}};
  GEN_116 = GEN_276[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_277 = {1{$random}};
  GEN_117 = GEN_277[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_278 = {1{$random}};
  GEN_118 = GEN_278[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_279 = {1{$random}};
  GEN_119 = GEN_279[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_280 = {1{$random}};
  GEN_120 = GEN_280[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_281 = {1{$random}};
  GEN_121 = GEN_281[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_282 = {1{$random}};
  GEN_122 = GEN_282[15:0];
  `endif
  `ifdef RANDOMIZE
  GEN_283 = {2{$random}};
  GEN_123 = GEN_283[37:0];
  `endif
  `ifdef RANDOMIZE
  GEN_284 = {1{$random}};
  GEN_124 = GEN_284[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_285 = {1{$random}};
  GEN_125 = GEN_285[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_286 = {1{$random}};
  GEN_126 = GEN_286[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_287 = {1{$random}};
  GEN_127 = GEN_287[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_288 = {1{$random}};
  GEN_128 = GEN_288[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_289 = {1{$random}};
  GEN_129 = GEN_289[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_290 = {1{$random}};
  GEN_130 = GEN_290[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_291 = {1{$random}};
  GEN_131 = GEN_291[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_292 = {1{$random}};
  GEN_132 = GEN_292[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_293 = {1{$random}};
  GEN_133 = GEN_293[6:0];
  `endif
  `ifdef RANDOMIZE
  GEN_294 = {1{$random}};
  GEN_134 = GEN_294[21:0];
  `endif
  `ifdef RANDOMIZE
  GEN_295 = {1{$random}};
  GEN_135 = GEN_295[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_296 = {1{$random}};
  GEN_136 = GEN_296[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_297 = {1{$random}};
  GEN_137 = GEN_297[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_298 = {1{$random}};
  GEN_138 = GEN_298[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_299 = {1{$random}};
  GEN_139 = GEN_299[30:0];
  `endif
  `ifdef RANDOMIZE
  GEN_300 = {1{$random}};
  GEN_140 = GEN_300[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_301 = {1{$random}};
  GEN_141 = GEN_301[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_302 = {1{$random}};
  GEN_142 = GEN_302[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_303 = {1{$random}};
  GEN_143 = GEN_303[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_304 = {1{$random}};
  GEN_144 = GEN_304[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_305 = {1{$random}};
  GEN_145 = GEN_305[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_306 = {1{$random}};
  GEN_146 = GEN_306[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_307 = {1{$random}};
  GEN_147 = GEN_307[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_308 = {1{$random}};
  GEN_148 = GEN_308[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_309 = {1{$random}};
  GEN_149 = GEN_309[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_310 = {1{$random}};
  GEN_150 = GEN_310[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_311 = {1{$random}};
  GEN_151 = GEN_311[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_312 = {1{$random}};
  GEN_152 = GEN_312[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_313 = {1{$random}};
  GEN_153 = GEN_313[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_314 = {1{$random}};
  GEN_154 = GEN_314[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_315 = {1{$random}};
  GEN_155 = GEN_315[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_316 = {1{$random}};
  GEN_156 = GEN_316[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_317 = {1{$random}};
  GEN_157 = GEN_317[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_318 = {1{$random}};
  GEN_158 = GEN_318[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_319 = {1{$random}};
  GEN_159 = GEN_319[0:0];
  `endif
  end
`endif
endmodule
module Queue(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_header_src,
  input  [1:0] io_enq_bits_header_dst,
  input  [25:0] io_enq_bits_payload_addr_block,
  input   io_enq_bits_payload_client_xact_id,
  input  [2:0] io_enq_bits_payload_addr_beat,
  input   io_enq_bits_payload_is_builtin_type,
  input  [2:0] io_enq_bits_payload_a_type,
  input  [11:0] io_enq_bits_payload_union,
  input  [63:0] io_enq_bits_payload_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_header_src,
  output [1:0] io_deq_bits_header_dst,
  output [25:0] io_deq_bits_payload_addr_block,
  output  io_deq_bits_payload_client_xact_id,
  output [2:0] io_deq_bits_payload_addr_beat,
  output  io_deq_bits_payload_is_builtin_type,
  output [2:0] io_deq_bits_payload_a_type,
  output [11:0] io_deq_bits_payload_union,
  output [63:0] io_deq_bits_payload_data,
  output  io_count
);
  reg [1:0] ram_header_src [0:0];
  reg [31:0] GEN_0;
  wire [1:0] ram_header_src_T_1144_data;
  wire  ram_header_src_T_1144_addr;
  wire  ram_header_src_T_1144_en;
  wire [1:0] ram_header_src_T_1025_data;
  wire  ram_header_src_T_1025_addr;
  wire  ram_header_src_T_1025_mask;
  wire  ram_header_src_T_1025_en;
  reg [1:0] ram_header_dst [0:0];
  reg [31:0] GEN_1;
  wire [1:0] ram_header_dst_T_1144_data;
  wire  ram_header_dst_T_1144_addr;
  wire  ram_header_dst_T_1144_en;
  wire [1:0] ram_header_dst_T_1025_data;
  wire  ram_header_dst_T_1025_addr;
  wire  ram_header_dst_T_1025_mask;
  wire  ram_header_dst_T_1025_en;
  reg [25:0] ram_payload_addr_block [0:0];
  reg [31:0] GEN_2;
  wire [25:0] ram_payload_addr_block_T_1144_data;
  wire  ram_payload_addr_block_T_1144_addr;
  wire  ram_payload_addr_block_T_1144_en;
  wire [25:0] ram_payload_addr_block_T_1025_data;
  wire  ram_payload_addr_block_T_1025_addr;
  wire  ram_payload_addr_block_T_1025_mask;
  wire  ram_payload_addr_block_T_1025_en;
  reg  ram_payload_client_xact_id [0:0];
  reg [31:0] GEN_3;
  wire  ram_payload_client_xact_id_T_1144_data;
  wire  ram_payload_client_xact_id_T_1144_addr;
  wire  ram_payload_client_xact_id_T_1144_en;
  wire  ram_payload_client_xact_id_T_1025_data;
  wire  ram_payload_client_xact_id_T_1025_addr;
  wire  ram_payload_client_xact_id_T_1025_mask;
  wire  ram_payload_client_xact_id_T_1025_en;
  reg [2:0] ram_payload_addr_beat [0:0];
  reg [31:0] GEN_4;
  wire [2:0] ram_payload_addr_beat_T_1144_data;
  wire  ram_payload_addr_beat_T_1144_addr;
  wire  ram_payload_addr_beat_T_1144_en;
  wire [2:0] ram_payload_addr_beat_T_1025_data;
  wire  ram_payload_addr_beat_T_1025_addr;
  wire  ram_payload_addr_beat_T_1025_mask;
  wire  ram_payload_addr_beat_T_1025_en;
  reg  ram_payload_is_builtin_type [0:0];
  reg [31:0] GEN_5;
  wire  ram_payload_is_builtin_type_T_1144_data;
  wire  ram_payload_is_builtin_type_T_1144_addr;
  wire  ram_payload_is_builtin_type_T_1144_en;
  wire  ram_payload_is_builtin_type_T_1025_data;
  wire  ram_payload_is_builtin_type_T_1025_addr;
  wire  ram_payload_is_builtin_type_T_1025_mask;
  wire  ram_payload_is_builtin_type_T_1025_en;
  reg [2:0] ram_payload_a_type [0:0];
  reg [31:0] GEN_6;
  wire [2:0] ram_payload_a_type_T_1144_data;
  wire  ram_payload_a_type_T_1144_addr;
  wire  ram_payload_a_type_T_1144_en;
  wire [2:0] ram_payload_a_type_T_1025_data;
  wire  ram_payload_a_type_T_1025_addr;
  wire  ram_payload_a_type_T_1025_mask;
  wire  ram_payload_a_type_T_1025_en;
  reg [11:0] ram_payload_union [0:0];
  reg [31:0] GEN_7;
  wire [11:0] ram_payload_union_T_1144_data;
  wire  ram_payload_union_T_1144_addr;
  wire  ram_payload_union_T_1144_en;
  wire [11:0] ram_payload_union_T_1025_data;
  wire  ram_payload_union_T_1025_addr;
  wire  ram_payload_union_T_1025_mask;
  wire  ram_payload_union_T_1025_en;
  reg [63:0] ram_payload_data [0:0];
  reg [63:0] GEN_8;
  wire [63:0] ram_payload_data_T_1144_data;
  wire  ram_payload_data_T_1144_addr;
  wire  ram_payload_data_T_1144_en;
  wire [63:0] ram_payload_data_T_1025_data;
  wire  ram_payload_data_T_1025_addr;
  wire  ram_payload_data_T_1025_mask;
  wire  ram_payload_data_T_1025_en;
  reg  maybe_full;
  reg [31:0] GEN_9;
  wire  T_1022;
  wire  T_1023;
  wire  do_enq;
  wire  T_1024;
  wire  do_deq;
  wire  T_1139;
  wire  GEN_21;
  wire  T_1141;
  wire [1:0] T_1256;
  wire  ptr_diff;
  wire [1:0] T_1258;
  assign io_enq_ready = T_1022;
  assign io_deq_valid = T_1141;
  assign io_deq_bits_header_src = ram_header_src_T_1144_data;
  assign io_deq_bits_header_dst = ram_header_dst_T_1144_data;
  assign io_deq_bits_payload_addr_block = ram_payload_addr_block_T_1144_data;
  assign io_deq_bits_payload_client_xact_id = ram_payload_client_xact_id_T_1144_data;
  assign io_deq_bits_payload_addr_beat = ram_payload_addr_beat_T_1144_data;
  assign io_deq_bits_payload_is_builtin_type = ram_payload_is_builtin_type_T_1144_data;
  assign io_deq_bits_payload_a_type = ram_payload_a_type_T_1144_data;
  assign io_deq_bits_payload_union = ram_payload_union_T_1144_data;
  assign io_deq_bits_payload_data = ram_payload_data_T_1144_data;
  assign io_count = T_1258[0];
  assign ram_header_src_T_1144_addr = 1'h0;
  assign ram_header_src_T_1144_en = 1'h1;
  assign ram_header_src_T_1144_data = ram_header_src[ram_header_src_T_1144_addr];
  assign ram_header_src_T_1025_data = io_enq_bits_header_src;
  assign ram_header_src_T_1025_addr = 1'h0;
  assign ram_header_src_T_1025_mask = do_enq;
  assign ram_header_src_T_1025_en = do_enq;
  assign ram_header_dst_T_1144_addr = 1'h0;
  assign ram_header_dst_T_1144_en = 1'h1;
  assign ram_header_dst_T_1144_data = ram_header_dst[ram_header_dst_T_1144_addr];
  assign ram_header_dst_T_1025_data = io_enq_bits_header_dst;
  assign ram_header_dst_T_1025_addr = 1'h0;
  assign ram_header_dst_T_1025_mask = do_enq;
  assign ram_header_dst_T_1025_en = do_enq;
  assign ram_payload_addr_block_T_1144_addr = 1'h0;
  assign ram_payload_addr_block_T_1144_en = 1'h1;
  assign ram_payload_addr_block_T_1144_data = ram_payload_addr_block[ram_payload_addr_block_T_1144_addr];
  assign ram_payload_addr_block_T_1025_data = io_enq_bits_payload_addr_block;
  assign ram_payload_addr_block_T_1025_addr = 1'h0;
  assign ram_payload_addr_block_T_1025_mask = do_enq;
  assign ram_payload_addr_block_T_1025_en = do_enq;
  assign ram_payload_client_xact_id_T_1144_addr = 1'h0;
  assign ram_payload_client_xact_id_T_1144_en = 1'h1;
  assign ram_payload_client_xact_id_T_1144_data = ram_payload_client_xact_id[ram_payload_client_xact_id_T_1144_addr];
  assign ram_payload_client_xact_id_T_1025_data = io_enq_bits_payload_client_xact_id;
  assign ram_payload_client_xact_id_T_1025_addr = 1'h0;
  assign ram_payload_client_xact_id_T_1025_mask = do_enq;
  assign ram_payload_client_xact_id_T_1025_en = do_enq;
  assign ram_payload_addr_beat_T_1144_addr = 1'h0;
  assign ram_payload_addr_beat_T_1144_en = 1'h1;
  assign ram_payload_addr_beat_T_1144_data = ram_payload_addr_beat[ram_payload_addr_beat_T_1144_addr];
  assign ram_payload_addr_beat_T_1025_data = io_enq_bits_payload_addr_beat;
  assign ram_payload_addr_beat_T_1025_addr = 1'h0;
  assign ram_payload_addr_beat_T_1025_mask = do_enq;
  assign ram_payload_addr_beat_T_1025_en = do_enq;
  assign ram_payload_is_builtin_type_T_1144_addr = 1'h0;
  assign ram_payload_is_builtin_type_T_1144_en = 1'h1;
  assign ram_payload_is_builtin_type_T_1144_data = ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1144_addr];
  assign ram_payload_is_builtin_type_T_1025_data = io_enq_bits_payload_is_builtin_type;
  assign ram_payload_is_builtin_type_T_1025_addr = 1'h0;
  assign ram_payload_is_builtin_type_T_1025_mask = do_enq;
  assign ram_payload_is_builtin_type_T_1025_en = do_enq;
  assign ram_payload_a_type_T_1144_addr = 1'h0;
  assign ram_payload_a_type_T_1144_en = 1'h1;
  assign ram_payload_a_type_T_1144_data = ram_payload_a_type[ram_payload_a_type_T_1144_addr];
  assign ram_payload_a_type_T_1025_data = io_enq_bits_payload_a_type;
  assign ram_payload_a_type_T_1025_addr = 1'h0;
  assign ram_payload_a_type_T_1025_mask = do_enq;
  assign ram_payload_a_type_T_1025_en = do_enq;
  assign ram_payload_union_T_1144_addr = 1'h0;
  assign ram_payload_union_T_1144_en = 1'h1;
  assign ram_payload_union_T_1144_data = ram_payload_union[ram_payload_union_T_1144_addr];
  assign ram_payload_union_T_1025_data = io_enq_bits_payload_union;
  assign ram_payload_union_T_1025_addr = 1'h0;
  assign ram_payload_union_T_1025_mask = do_enq;
  assign ram_payload_union_T_1025_en = do_enq;
  assign ram_payload_data_T_1144_addr = 1'h0;
  assign ram_payload_data_T_1144_en = 1'h1;
  assign ram_payload_data_T_1144_data = ram_payload_data[ram_payload_data_T_1144_addr];
  assign ram_payload_data_T_1025_data = io_enq_bits_payload_data;
  assign ram_payload_data_T_1025_addr = 1'h0;
  assign ram_payload_data_T_1025_mask = do_enq;
  assign ram_payload_data_T_1025_en = do_enq;
  assign T_1022 = maybe_full == 1'h0;
  assign T_1023 = io_enq_ready & io_enq_valid;
  assign do_enq = T_1023;
  assign T_1024 = io_deq_ready & io_deq_valid;
  assign do_deq = T_1024;
  assign T_1139 = do_enq != do_deq;
  assign GEN_21 = T_1139 ? do_enq : maybe_full;
  assign T_1141 = T_1022 == 1'h0;
  assign T_1256 = 1'h0 - 1'h0;
  assign ptr_diff = T_1256[0:0];
  assign T_1258 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_header_src[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_header_dst[initvar] = GEN_1[1:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_addr_block[initvar] = GEN_2[25:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_client_xact_id[initvar] = GEN_3[0:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_addr_beat[initvar] = GEN_4[2:0];
  `endif
  GEN_5 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_is_builtin_type[initvar] = GEN_5[0:0];
  `endif
  GEN_6 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_a_type[initvar] = GEN_6[2:0];
  `endif
  GEN_7 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_union[initvar] = GEN_7[11:0];
  `endif
  GEN_8 = {2{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_data[initvar] = GEN_8[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_9 = {1{$random}};
  maybe_full = GEN_9[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_header_src_T_1025_en & ram_header_src_T_1025_mask) begin
      ram_header_src[ram_header_src_T_1025_addr] <= ram_header_src_T_1025_data;
    end
    if(ram_header_dst_T_1025_en & ram_header_dst_T_1025_mask) begin
      ram_header_dst[ram_header_dst_T_1025_addr] <= ram_header_dst_T_1025_data;
    end
    if(ram_payload_addr_block_T_1025_en & ram_payload_addr_block_T_1025_mask) begin
      ram_payload_addr_block[ram_payload_addr_block_T_1025_addr] <= ram_payload_addr_block_T_1025_data;
    end
    if(ram_payload_client_xact_id_T_1025_en & ram_payload_client_xact_id_T_1025_mask) begin
      ram_payload_client_xact_id[ram_payload_client_xact_id_T_1025_addr] <= ram_payload_client_xact_id_T_1025_data;
    end
    if(ram_payload_addr_beat_T_1025_en & ram_payload_addr_beat_T_1025_mask) begin
      ram_payload_addr_beat[ram_payload_addr_beat_T_1025_addr] <= ram_payload_addr_beat_T_1025_data;
    end
    if(ram_payload_is_builtin_type_T_1025_en & ram_payload_is_builtin_type_T_1025_mask) begin
      ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1025_addr] <= ram_payload_is_builtin_type_T_1025_data;
    end
    if(ram_payload_a_type_T_1025_en & ram_payload_a_type_T_1025_mask) begin
      ram_payload_a_type[ram_payload_a_type_T_1025_addr] <= ram_payload_a_type_T_1025_data;
    end
    if(ram_payload_union_T_1025_en & ram_payload_union_T_1025_mask) begin
      ram_payload_union[ram_payload_union_T_1025_addr] <= ram_payload_union_T_1025_data;
    end
    if(ram_payload_data_T_1025_en & ram_payload_data_T_1025_mask) begin
      ram_payload_data[ram_payload_data_T_1025_addr] <= ram_payload_data_T_1025_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_1139) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_1(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_header_src,
  input  [1:0] io_enq_bits_header_dst,
  input  [25:0] io_enq_bits_payload_addr_block,
  input  [1:0] io_enq_bits_payload_p_type,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_header_src,
  output [1:0] io_deq_bits_header_dst,
  output [25:0] io_deq_bits_payload_addr_block,
  output [1:0] io_deq_bits_payload_p_type,
  output  io_count
);
  reg [1:0] ram_header_src [0:0];
  reg [31:0] GEN_0;
  wire [1:0] ram_header_src_T_1094_data;
  wire  ram_header_src_T_1094_addr;
  wire  ram_header_src_T_1094_en;
  wire [1:0] ram_header_src_T_980_data;
  wire  ram_header_src_T_980_addr;
  wire  ram_header_src_T_980_mask;
  wire  ram_header_src_T_980_en;
  reg [1:0] ram_header_dst [0:0];
  reg [31:0] GEN_1;
  wire [1:0] ram_header_dst_T_1094_data;
  wire  ram_header_dst_T_1094_addr;
  wire  ram_header_dst_T_1094_en;
  wire [1:0] ram_header_dst_T_980_data;
  wire  ram_header_dst_T_980_addr;
  wire  ram_header_dst_T_980_mask;
  wire  ram_header_dst_T_980_en;
  reg [25:0] ram_payload_addr_block [0:0];
  reg [31:0] GEN_2;
  wire [25:0] ram_payload_addr_block_T_1094_data;
  wire  ram_payload_addr_block_T_1094_addr;
  wire  ram_payload_addr_block_T_1094_en;
  wire [25:0] ram_payload_addr_block_T_980_data;
  wire  ram_payload_addr_block_T_980_addr;
  wire  ram_payload_addr_block_T_980_mask;
  wire  ram_payload_addr_block_T_980_en;
  reg [1:0] ram_payload_p_type [0:0];
  reg [31:0] GEN_3;
  wire [1:0] ram_payload_p_type_T_1094_data;
  wire  ram_payload_p_type_T_1094_addr;
  wire  ram_payload_p_type_T_1094_en;
  wire [1:0] ram_payload_p_type_T_980_data;
  wire  ram_payload_p_type_T_980_addr;
  wire  ram_payload_p_type_T_980_mask;
  wire  ram_payload_p_type_T_980_en;
  reg  maybe_full;
  reg [31:0] GEN_4;
  wire  T_977;
  wire  T_978;
  wire  do_enq;
  wire  T_979;
  wire  do_deq;
  wire  T_1089;
  wire  GEN_11;
  wire  T_1091;
  wire [1:0] T_1201;
  wire  ptr_diff;
  wire [1:0] T_1203;
  assign io_enq_ready = T_977;
  assign io_deq_valid = T_1091;
  assign io_deq_bits_header_src = ram_header_src_T_1094_data;
  assign io_deq_bits_header_dst = ram_header_dst_T_1094_data;
  assign io_deq_bits_payload_addr_block = ram_payload_addr_block_T_1094_data;
  assign io_deq_bits_payload_p_type = ram_payload_p_type_T_1094_data;
  assign io_count = T_1203[0];
  assign ram_header_src_T_1094_addr = 1'h0;
  assign ram_header_src_T_1094_en = 1'h1;
  assign ram_header_src_T_1094_data = ram_header_src[ram_header_src_T_1094_addr];
  assign ram_header_src_T_980_data = io_enq_bits_header_src;
  assign ram_header_src_T_980_addr = 1'h0;
  assign ram_header_src_T_980_mask = do_enq;
  assign ram_header_src_T_980_en = do_enq;
  assign ram_header_dst_T_1094_addr = 1'h0;
  assign ram_header_dst_T_1094_en = 1'h1;
  assign ram_header_dst_T_1094_data = ram_header_dst[ram_header_dst_T_1094_addr];
  assign ram_header_dst_T_980_data = io_enq_bits_header_dst;
  assign ram_header_dst_T_980_addr = 1'h0;
  assign ram_header_dst_T_980_mask = do_enq;
  assign ram_header_dst_T_980_en = do_enq;
  assign ram_payload_addr_block_T_1094_addr = 1'h0;
  assign ram_payload_addr_block_T_1094_en = 1'h1;
  assign ram_payload_addr_block_T_1094_data = ram_payload_addr_block[ram_payload_addr_block_T_1094_addr];
  assign ram_payload_addr_block_T_980_data = io_enq_bits_payload_addr_block;
  assign ram_payload_addr_block_T_980_addr = 1'h0;
  assign ram_payload_addr_block_T_980_mask = do_enq;
  assign ram_payload_addr_block_T_980_en = do_enq;
  assign ram_payload_p_type_T_1094_addr = 1'h0;
  assign ram_payload_p_type_T_1094_en = 1'h1;
  assign ram_payload_p_type_T_1094_data = ram_payload_p_type[ram_payload_p_type_T_1094_addr];
  assign ram_payload_p_type_T_980_data = io_enq_bits_payload_p_type;
  assign ram_payload_p_type_T_980_addr = 1'h0;
  assign ram_payload_p_type_T_980_mask = do_enq;
  assign ram_payload_p_type_T_980_en = do_enq;
  assign T_977 = maybe_full == 1'h0;
  assign T_978 = io_enq_ready & io_enq_valid;
  assign do_enq = T_978;
  assign T_979 = io_deq_ready & io_deq_valid;
  assign do_deq = T_979;
  assign T_1089 = do_enq != do_deq;
  assign GEN_11 = T_1089 ? do_enq : maybe_full;
  assign T_1091 = T_977 == 1'h0;
  assign T_1201 = 1'h0 - 1'h0;
  assign ptr_diff = T_1201[0:0];
  assign T_1203 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_header_src[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_header_dst[initvar] = GEN_1[1:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_addr_block[initvar] = GEN_2[25:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_p_type[initvar] = GEN_3[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_4 = {1{$random}};
  maybe_full = GEN_4[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_header_src_T_980_en & ram_header_src_T_980_mask) begin
      ram_header_src[ram_header_src_T_980_addr] <= ram_header_src_T_980_data;
    end
    if(ram_header_dst_T_980_en & ram_header_dst_T_980_mask) begin
      ram_header_dst[ram_header_dst_T_980_addr] <= ram_header_dst_T_980_data;
    end
    if(ram_payload_addr_block_T_980_en & ram_payload_addr_block_T_980_mask) begin
      ram_payload_addr_block[ram_payload_addr_block_T_980_addr] <= ram_payload_addr_block_T_980_data;
    end
    if(ram_payload_p_type_T_980_en & ram_payload_p_type_T_980_mask) begin
      ram_payload_p_type[ram_payload_p_type_T_980_addr] <= ram_payload_p_type_T_980_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_1089) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_2(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_header_src,
  input  [1:0] io_enq_bits_header_dst,
  input  [2:0] io_enq_bits_payload_addr_beat,
  input  [25:0] io_enq_bits_payload_addr_block,
  input   io_enq_bits_payload_client_xact_id,
  input   io_enq_bits_payload_voluntary,
  input  [2:0] io_enq_bits_payload_r_type,
  input  [63:0] io_enq_bits_payload_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_header_src,
  output [1:0] io_deq_bits_header_dst,
  output [2:0] io_deq_bits_payload_addr_beat,
  output [25:0] io_deq_bits_payload_addr_block,
  output  io_deq_bits_payload_client_xact_id,
  output  io_deq_bits_payload_voluntary,
  output [2:0] io_deq_bits_payload_r_type,
  output [63:0] io_deq_bits_payload_data,
  output [1:0] io_count
);
  reg [1:0] ram_header_src [0:1];
  reg [31:0] GEN_0;
  wire [1:0] ram_header_src_T_1144_data;
  wire  ram_header_src_T_1144_addr;
  wire  ram_header_src_T_1144_en;
  wire [1:0] ram_header_src_T_1018_data;
  wire  ram_header_src_T_1018_addr;
  wire  ram_header_src_T_1018_mask;
  wire  ram_header_src_T_1018_en;
  reg [1:0] ram_header_dst [0:1];
  reg [31:0] GEN_1;
  wire [1:0] ram_header_dst_T_1144_data;
  wire  ram_header_dst_T_1144_addr;
  wire  ram_header_dst_T_1144_en;
  wire [1:0] ram_header_dst_T_1018_data;
  wire  ram_header_dst_T_1018_addr;
  wire  ram_header_dst_T_1018_mask;
  wire  ram_header_dst_T_1018_en;
  reg [2:0] ram_payload_addr_beat [0:1];
  reg [31:0] GEN_2;
  wire [2:0] ram_payload_addr_beat_T_1144_data;
  wire  ram_payload_addr_beat_T_1144_addr;
  wire  ram_payload_addr_beat_T_1144_en;
  wire [2:0] ram_payload_addr_beat_T_1018_data;
  wire  ram_payload_addr_beat_T_1018_addr;
  wire  ram_payload_addr_beat_T_1018_mask;
  wire  ram_payload_addr_beat_T_1018_en;
  reg [25:0] ram_payload_addr_block [0:1];
  reg [31:0] GEN_3;
  wire [25:0] ram_payload_addr_block_T_1144_data;
  wire  ram_payload_addr_block_T_1144_addr;
  wire  ram_payload_addr_block_T_1144_en;
  wire [25:0] ram_payload_addr_block_T_1018_data;
  wire  ram_payload_addr_block_T_1018_addr;
  wire  ram_payload_addr_block_T_1018_mask;
  wire  ram_payload_addr_block_T_1018_en;
  reg  ram_payload_client_xact_id [0:1];
  reg [31:0] GEN_4;
  wire  ram_payload_client_xact_id_T_1144_data;
  wire  ram_payload_client_xact_id_T_1144_addr;
  wire  ram_payload_client_xact_id_T_1144_en;
  wire  ram_payload_client_xact_id_T_1018_data;
  wire  ram_payload_client_xact_id_T_1018_addr;
  wire  ram_payload_client_xact_id_T_1018_mask;
  wire  ram_payload_client_xact_id_T_1018_en;
  reg  ram_payload_voluntary [0:1];
  reg [31:0] GEN_5;
  wire  ram_payload_voluntary_T_1144_data;
  wire  ram_payload_voluntary_T_1144_addr;
  wire  ram_payload_voluntary_T_1144_en;
  wire  ram_payload_voluntary_T_1018_data;
  wire  ram_payload_voluntary_T_1018_addr;
  wire  ram_payload_voluntary_T_1018_mask;
  wire  ram_payload_voluntary_T_1018_en;
  reg [2:0] ram_payload_r_type [0:1];
  reg [31:0] GEN_6;
  wire [2:0] ram_payload_r_type_T_1144_data;
  wire  ram_payload_r_type_T_1144_addr;
  wire  ram_payload_r_type_T_1144_en;
  wire [2:0] ram_payload_r_type_T_1018_data;
  wire  ram_payload_r_type_T_1018_addr;
  wire  ram_payload_r_type_T_1018_mask;
  wire  ram_payload_r_type_T_1018_en;
  reg [63:0] ram_payload_data [0:1];
  reg [63:0] GEN_7;
  wire [63:0] ram_payload_data_T_1144_data;
  wire  ram_payload_data_T_1144_addr;
  wire  ram_payload_data_T_1144_en;
  wire [63:0] ram_payload_data_T_1018_data;
  wire  ram_payload_data_T_1018_addr;
  wire  ram_payload_data_T_1018_mask;
  wire  ram_payload_data_T_1018_en;
  reg  T_1010;
  reg [31:0] GEN_8;
  reg  T_1012;
  reg [31:0] GEN_9;
  reg  maybe_full;
  reg [31:0] GEN_10;
  wire  ptr_match;
  wire  T_1015;
  wire  empty;
  wire  full;
  wire  T_1016;
  wire  do_enq;
  wire  T_1017;
  wire  do_deq;
  wire [1:0] T_1132;
  wire  T_1133;
  wire  GEN_19;
  wire [1:0] T_1137;
  wire  T_1138;
  wire  GEN_20;
  wire  T_1139;
  wire  GEN_21;
  wire  T_1141;
  wire  T_1143;
  wire [1:0] T_1255;
  wire  ptr_diff;
  wire  T_1256;
  wire [1:0] T_1257;
  assign io_enq_ready = T_1143;
  assign io_deq_valid = T_1141;
  assign io_deq_bits_header_src = ram_header_src_T_1144_data;
  assign io_deq_bits_header_dst = ram_header_dst_T_1144_data;
  assign io_deq_bits_payload_addr_beat = ram_payload_addr_beat_T_1144_data;
  assign io_deq_bits_payload_addr_block = ram_payload_addr_block_T_1144_data;
  assign io_deq_bits_payload_client_xact_id = ram_payload_client_xact_id_T_1144_data;
  assign io_deq_bits_payload_voluntary = ram_payload_voluntary_T_1144_data;
  assign io_deq_bits_payload_r_type = ram_payload_r_type_T_1144_data;
  assign io_deq_bits_payload_data = ram_payload_data_T_1144_data;
  assign io_count = T_1257;
  assign ram_header_src_T_1144_addr = T_1012;
  assign ram_header_src_T_1144_en = 1'h1;
  assign ram_header_src_T_1144_data = ram_header_src[ram_header_src_T_1144_addr];
  assign ram_header_src_T_1018_data = io_enq_bits_header_src;
  assign ram_header_src_T_1018_addr = T_1010;
  assign ram_header_src_T_1018_mask = do_enq;
  assign ram_header_src_T_1018_en = do_enq;
  assign ram_header_dst_T_1144_addr = T_1012;
  assign ram_header_dst_T_1144_en = 1'h1;
  assign ram_header_dst_T_1144_data = ram_header_dst[ram_header_dst_T_1144_addr];
  assign ram_header_dst_T_1018_data = io_enq_bits_header_dst;
  assign ram_header_dst_T_1018_addr = T_1010;
  assign ram_header_dst_T_1018_mask = do_enq;
  assign ram_header_dst_T_1018_en = do_enq;
  assign ram_payload_addr_beat_T_1144_addr = T_1012;
  assign ram_payload_addr_beat_T_1144_en = 1'h1;
  assign ram_payload_addr_beat_T_1144_data = ram_payload_addr_beat[ram_payload_addr_beat_T_1144_addr];
  assign ram_payload_addr_beat_T_1018_data = io_enq_bits_payload_addr_beat;
  assign ram_payload_addr_beat_T_1018_addr = T_1010;
  assign ram_payload_addr_beat_T_1018_mask = do_enq;
  assign ram_payload_addr_beat_T_1018_en = do_enq;
  assign ram_payload_addr_block_T_1144_addr = T_1012;
  assign ram_payload_addr_block_T_1144_en = 1'h1;
  assign ram_payload_addr_block_T_1144_data = ram_payload_addr_block[ram_payload_addr_block_T_1144_addr];
  assign ram_payload_addr_block_T_1018_data = io_enq_bits_payload_addr_block;
  assign ram_payload_addr_block_T_1018_addr = T_1010;
  assign ram_payload_addr_block_T_1018_mask = do_enq;
  assign ram_payload_addr_block_T_1018_en = do_enq;
  assign ram_payload_client_xact_id_T_1144_addr = T_1012;
  assign ram_payload_client_xact_id_T_1144_en = 1'h1;
  assign ram_payload_client_xact_id_T_1144_data = ram_payload_client_xact_id[ram_payload_client_xact_id_T_1144_addr];
  assign ram_payload_client_xact_id_T_1018_data = io_enq_bits_payload_client_xact_id;
  assign ram_payload_client_xact_id_T_1018_addr = T_1010;
  assign ram_payload_client_xact_id_T_1018_mask = do_enq;
  assign ram_payload_client_xact_id_T_1018_en = do_enq;
  assign ram_payload_voluntary_T_1144_addr = T_1012;
  assign ram_payload_voluntary_T_1144_en = 1'h1;
  assign ram_payload_voluntary_T_1144_data = ram_payload_voluntary[ram_payload_voluntary_T_1144_addr];
  assign ram_payload_voluntary_T_1018_data = io_enq_bits_payload_voluntary;
  assign ram_payload_voluntary_T_1018_addr = T_1010;
  assign ram_payload_voluntary_T_1018_mask = do_enq;
  assign ram_payload_voluntary_T_1018_en = do_enq;
  assign ram_payload_r_type_T_1144_addr = T_1012;
  assign ram_payload_r_type_T_1144_en = 1'h1;
  assign ram_payload_r_type_T_1144_data = ram_payload_r_type[ram_payload_r_type_T_1144_addr];
  assign ram_payload_r_type_T_1018_data = io_enq_bits_payload_r_type;
  assign ram_payload_r_type_T_1018_addr = T_1010;
  assign ram_payload_r_type_T_1018_mask = do_enq;
  assign ram_payload_r_type_T_1018_en = do_enq;
  assign ram_payload_data_T_1144_addr = T_1012;
  assign ram_payload_data_T_1144_en = 1'h1;
  assign ram_payload_data_T_1144_data = ram_payload_data[ram_payload_data_T_1144_addr];
  assign ram_payload_data_T_1018_data = io_enq_bits_payload_data;
  assign ram_payload_data_T_1018_addr = T_1010;
  assign ram_payload_data_T_1018_mask = do_enq;
  assign ram_payload_data_T_1018_en = do_enq;
  assign ptr_match = T_1010 == T_1012;
  assign T_1015 = maybe_full == 1'h0;
  assign empty = ptr_match & T_1015;
  assign full = ptr_match & maybe_full;
  assign T_1016 = io_enq_ready & io_enq_valid;
  assign do_enq = T_1016;
  assign T_1017 = io_deq_ready & io_deq_valid;
  assign do_deq = T_1017;
  assign T_1132 = T_1010 + 1'h1;
  assign T_1133 = T_1132[0:0];
  assign GEN_19 = do_enq ? T_1133 : T_1010;
  assign T_1137 = T_1012 + 1'h1;
  assign T_1138 = T_1137[0:0];
  assign GEN_20 = do_deq ? T_1138 : T_1012;
  assign T_1139 = do_enq != do_deq;
  assign GEN_21 = T_1139 ? do_enq : maybe_full;
  assign T_1141 = empty == 1'h0;
  assign T_1143 = full == 1'h0;
  assign T_1255 = T_1010 - T_1012;
  assign ptr_diff = T_1255[0:0];
  assign T_1256 = maybe_full & ptr_match;
  assign T_1257 = {T_1256,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_header_src[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_header_dst[initvar] = GEN_1[1:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_addr_beat[initvar] = GEN_2[2:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_addr_block[initvar] = GEN_3[25:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_client_xact_id[initvar] = GEN_4[0:0];
  `endif
  GEN_5 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_voluntary[initvar] = GEN_5[0:0];
  `endif
  GEN_6 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_r_type[initvar] = GEN_6[2:0];
  `endif
  GEN_7 = {2{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_data[initvar] = GEN_7[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_8 = {1{$random}};
  T_1010 = GEN_8[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_9 = {1{$random}};
  T_1012 = GEN_9[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_10 = {1{$random}};
  maybe_full = GEN_10[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_header_src_T_1018_en & ram_header_src_T_1018_mask) begin
      ram_header_src[ram_header_src_T_1018_addr] <= ram_header_src_T_1018_data;
    end
    if(ram_header_dst_T_1018_en & ram_header_dst_T_1018_mask) begin
      ram_header_dst[ram_header_dst_T_1018_addr] <= ram_header_dst_T_1018_data;
    end
    if(ram_payload_addr_beat_T_1018_en & ram_payload_addr_beat_T_1018_mask) begin
      ram_payload_addr_beat[ram_payload_addr_beat_T_1018_addr] <= ram_payload_addr_beat_T_1018_data;
    end
    if(ram_payload_addr_block_T_1018_en & ram_payload_addr_block_T_1018_mask) begin
      ram_payload_addr_block[ram_payload_addr_block_T_1018_addr] <= ram_payload_addr_block_T_1018_data;
    end
    if(ram_payload_client_xact_id_T_1018_en & ram_payload_client_xact_id_T_1018_mask) begin
      ram_payload_client_xact_id[ram_payload_client_xact_id_T_1018_addr] <= ram_payload_client_xact_id_T_1018_data;
    end
    if(ram_payload_voluntary_T_1018_en & ram_payload_voluntary_T_1018_mask) begin
      ram_payload_voluntary[ram_payload_voluntary_T_1018_addr] <= ram_payload_voluntary_T_1018_data;
    end
    if(ram_payload_r_type_T_1018_en & ram_payload_r_type_T_1018_mask) begin
      ram_payload_r_type[ram_payload_r_type_T_1018_addr] <= ram_payload_r_type_T_1018_data;
    end
    if(ram_payload_data_T_1018_en & ram_payload_data_T_1018_mask) begin
      ram_payload_data[ram_payload_data_T_1018_addr] <= ram_payload_data_T_1018_data;
    end
    if(reset) begin
      T_1010 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_1010 <= T_1133;
      end
    end
    if(reset) begin
      T_1012 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_1012 <= T_1138;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_1139) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_3(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_header_src,
  input  [1:0] io_enq_bits_header_dst,
  input  [2:0] io_enq_bits_payload_addr_beat,
  input   io_enq_bits_payload_client_xact_id,
  input  [1:0] io_enq_bits_payload_manager_xact_id,
  input   io_enq_bits_payload_is_builtin_type,
  input  [3:0] io_enq_bits_payload_g_type,
  input  [63:0] io_enq_bits_payload_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_header_src,
  output [1:0] io_deq_bits_header_dst,
  output [2:0] io_deq_bits_payload_addr_beat,
  output  io_deq_bits_payload_client_xact_id,
  output [1:0] io_deq_bits_payload_manager_xact_id,
  output  io_deq_bits_payload_is_builtin_type,
  output [3:0] io_deq_bits_payload_g_type,
  output [63:0] io_deq_bits_payload_data,
  output [1:0] io_count
);
  reg [1:0] ram_header_src [0:1];
  reg [31:0] GEN_0;
  wire [1:0] ram_header_src_T_1144_data;
  wire  ram_header_src_T_1144_addr;
  wire  ram_header_src_T_1144_en;
  wire [1:0] ram_header_src_T_1018_data;
  wire  ram_header_src_T_1018_addr;
  wire  ram_header_src_T_1018_mask;
  wire  ram_header_src_T_1018_en;
  reg [1:0] ram_header_dst [0:1];
  reg [31:0] GEN_1;
  wire [1:0] ram_header_dst_T_1144_data;
  wire  ram_header_dst_T_1144_addr;
  wire  ram_header_dst_T_1144_en;
  wire [1:0] ram_header_dst_T_1018_data;
  wire  ram_header_dst_T_1018_addr;
  wire  ram_header_dst_T_1018_mask;
  wire  ram_header_dst_T_1018_en;
  reg [2:0] ram_payload_addr_beat [0:1];
  reg [31:0] GEN_2;
  wire [2:0] ram_payload_addr_beat_T_1144_data;
  wire  ram_payload_addr_beat_T_1144_addr;
  wire  ram_payload_addr_beat_T_1144_en;
  wire [2:0] ram_payload_addr_beat_T_1018_data;
  wire  ram_payload_addr_beat_T_1018_addr;
  wire  ram_payload_addr_beat_T_1018_mask;
  wire  ram_payload_addr_beat_T_1018_en;
  reg  ram_payload_client_xact_id [0:1];
  reg [31:0] GEN_3;
  wire  ram_payload_client_xact_id_T_1144_data;
  wire  ram_payload_client_xact_id_T_1144_addr;
  wire  ram_payload_client_xact_id_T_1144_en;
  wire  ram_payload_client_xact_id_T_1018_data;
  wire  ram_payload_client_xact_id_T_1018_addr;
  wire  ram_payload_client_xact_id_T_1018_mask;
  wire  ram_payload_client_xact_id_T_1018_en;
  reg [1:0] ram_payload_manager_xact_id [0:1];
  reg [31:0] GEN_4;
  wire [1:0] ram_payload_manager_xact_id_T_1144_data;
  wire  ram_payload_manager_xact_id_T_1144_addr;
  wire  ram_payload_manager_xact_id_T_1144_en;
  wire [1:0] ram_payload_manager_xact_id_T_1018_data;
  wire  ram_payload_manager_xact_id_T_1018_addr;
  wire  ram_payload_manager_xact_id_T_1018_mask;
  wire  ram_payload_manager_xact_id_T_1018_en;
  reg  ram_payload_is_builtin_type [0:1];
  reg [31:0] GEN_5;
  wire  ram_payload_is_builtin_type_T_1144_data;
  wire  ram_payload_is_builtin_type_T_1144_addr;
  wire  ram_payload_is_builtin_type_T_1144_en;
  wire  ram_payload_is_builtin_type_T_1018_data;
  wire  ram_payload_is_builtin_type_T_1018_addr;
  wire  ram_payload_is_builtin_type_T_1018_mask;
  wire  ram_payload_is_builtin_type_T_1018_en;
  reg [3:0] ram_payload_g_type [0:1];
  reg [31:0] GEN_6;
  wire [3:0] ram_payload_g_type_T_1144_data;
  wire  ram_payload_g_type_T_1144_addr;
  wire  ram_payload_g_type_T_1144_en;
  wire [3:0] ram_payload_g_type_T_1018_data;
  wire  ram_payload_g_type_T_1018_addr;
  wire  ram_payload_g_type_T_1018_mask;
  wire  ram_payload_g_type_T_1018_en;
  reg [63:0] ram_payload_data [0:1];
  reg [63:0] GEN_7;
  wire [63:0] ram_payload_data_T_1144_data;
  wire  ram_payload_data_T_1144_addr;
  wire  ram_payload_data_T_1144_en;
  wire [63:0] ram_payload_data_T_1018_data;
  wire  ram_payload_data_T_1018_addr;
  wire  ram_payload_data_T_1018_mask;
  wire  ram_payload_data_T_1018_en;
  reg  T_1010;
  reg [31:0] GEN_8;
  reg  T_1012;
  reg [31:0] GEN_9;
  reg  maybe_full;
  reg [31:0] GEN_10;
  wire  ptr_match;
  wire  T_1015;
  wire  empty;
  wire  full;
  wire  T_1016;
  wire  do_enq;
  wire  T_1017;
  wire  do_deq;
  wire [1:0] T_1132;
  wire  T_1133;
  wire  GEN_19;
  wire [1:0] T_1137;
  wire  T_1138;
  wire  GEN_20;
  wire  T_1139;
  wire  GEN_21;
  wire  T_1141;
  wire  T_1143;
  wire [1:0] T_1255;
  wire  ptr_diff;
  wire  T_1256;
  wire [1:0] T_1257;
  assign io_enq_ready = T_1143;
  assign io_deq_valid = T_1141;
  assign io_deq_bits_header_src = ram_header_src_T_1144_data;
  assign io_deq_bits_header_dst = ram_header_dst_T_1144_data;
  assign io_deq_bits_payload_addr_beat = ram_payload_addr_beat_T_1144_data;
  assign io_deq_bits_payload_client_xact_id = ram_payload_client_xact_id_T_1144_data;
  assign io_deq_bits_payload_manager_xact_id = ram_payload_manager_xact_id_T_1144_data;
  assign io_deq_bits_payload_is_builtin_type = ram_payload_is_builtin_type_T_1144_data;
  assign io_deq_bits_payload_g_type = ram_payload_g_type_T_1144_data;
  assign io_deq_bits_payload_data = ram_payload_data_T_1144_data;
  assign io_count = T_1257;
  assign ram_header_src_T_1144_addr = T_1012;
  assign ram_header_src_T_1144_en = 1'h1;
  assign ram_header_src_T_1144_data = ram_header_src[ram_header_src_T_1144_addr];
  assign ram_header_src_T_1018_data = io_enq_bits_header_src;
  assign ram_header_src_T_1018_addr = T_1010;
  assign ram_header_src_T_1018_mask = do_enq;
  assign ram_header_src_T_1018_en = do_enq;
  assign ram_header_dst_T_1144_addr = T_1012;
  assign ram_header_dst_T_1144_en = 1'h1;
  assign ram_header_dst_T_1144_data = ram_header_dst[ram_header_dst_T_1144_addr];
  assign ram_header_dst_T_1018_data = io_enq_bits_header_dst;
  assign ram_header_dst_T_1018_addr = T_1010;
  assign ram_header_dst_T_1018_mask = do_enq;
  assign ram_header_dst_T_1018_en = do_enq;
  assign ram_payload_addr_beat_T_1144_addr = T_1012;
  assign ram_payload_addr_beat_T_1144_en = 1'h1;
  assign ram_payload_addr_beat_T_1144_data = ram_payload_addr_beat[ram_payload_addr_beat_T_1144_addr];
  assign ram_payload_addr_beat_T_1018_data = io_enq_bits_payload_addr_beat;
  assign ram_payload_addr_beat_T_1018_addr = T_1010;
  assign ram_payload_addr_beat_T_1018_mask = do_enq;
  assign ram_payload_addr_beat_T_1018_en = do_enq;
  assign ram_payload_client_xact_id_T_1144_addr = T_1012;
  assign ram_payload_client_xact_id_T_1144_en = 1'h1;
  assign ram_payload_client_xact_id_T_1144_data = ram_payload_client_xact_id[ram_payload_client_xact_id_T_1144_addr];
  assign ram_payload_client_xact_id_T_1018_data = io_enq_bits_payload_client_xact_id;
  assign ram_payload_client_xact_id_T_1018_addr = T_1010;
  assign ram_payload_client_xact_id_T_1018_mask = do_enq;
  assign ram_payload_client_xact_id_T_1018_en = do_enq;
  assign ram_payload_manager_xact_id_T_1144_addr = T_1012;
  assign ram_payload_manager_xact_id_T_1144_en = 1'h1;
  assign ram_payload_manager_xact_id_T_1144_data = ram_payload_manager_xact_id[ram_payload_manager_xact_id_T_1144_addr];
  assign ram_payload_manager_xact_id_T_1018_data = io_enq_bits_payload_manager_xact_id;
  assign ram_payload_manager_xact_id_T_1018_addr = T_1010;
  assign ram_payload_manager_xact_id_T_1018_mask = do_enq;
  assign ram_payload_manager_xact_id_T_1018_en = do_enq;
  assign ram_payload_is_builtin_type_T_1144_addr = T_1012;
  assign ram_payload_is_builtin_type_T_1144_en = 1'h1;
  assign ram_payload_is_builtin_type_T_1144_data = ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1144_addr];
  assign ram_payload_is_builtin_type_T_1018_data = io_enq_bits_payload_is_builtin_type;
  assign ram_payload_is_builtin_type_T_1018_addr = T_1010;
  assign ram_payload_is_builtin_type_T_1018_mask = do_enq;
  assign ram_payload_is_builtin_type_T_1018_en = do_enq;
  assign ram_payload_g_type_T_1144_addr = T_1012;
  assign ram_payload_g_type_T_1144_en = 1'h1;
  assign ram_payload_g_type_T_1144_data = ram_payload_g_type[ram_payload_g_type_T_1144_addr];
  assign ram_payload_g_type_T_1018_data = io_enq_bits_payload_g_type;
  assign ram_payload_g_type_T_1018_addr = T_1010;
  assign ram_payload_g_type_T_1018_mask = do_enq;
  assign ram_payload_g_type_T_1018_en = do_enq;
  assign ram_payload_data_T_1144_addr = T_1012;
  assign ram_payload_data_T_1144_en = 1'h1;
  assign ram_payload_data_T_1144_data = ram_payload_data[ram_payload_data_T_1144_addr];
  assign ram_payload_data_T_1018_data = io_enq_bits_payload_data;
  assign ram_payload_data_T_1018_addr = T_1010;
  assign ram_payload_data_T_1018_mask = do_enq;
  assign ram_payload_data_T_1018_en = do_enq;
  assign ptr_match = T_1010 == T_1012;
  assign T_1015 = maybe_full == 1'h0;
  assign empty = ptr_match & T_1015;
  assign full = ptr_match & maybe_full;
  assign T_1016 = io_enq_ready & io_enq_valid;
  assign do_enq = T_1016;
  assign T_1017 = io_deq_ready & io_deq_valid;
  assign do_deq = T_1017;
  assign T_1132 = T_1010 + 1'h1;
  assign T_1133 = T_1132[0:0];
  assign GEN_19 = do_enq ? T_1133 : T_1010;
  assign T_1137 = T_1012 + 1'h1;
  assign T_1138 = T_1137[0:0];
  assign GEN_20 = do_deq ? T_1138 : T_1012;
  assign T_1139 = do_enq != do_deq;
  assign GEN_21 = T_1139 ? do_enq : maybe_full;
  assign T_1141 = empty == 1'h0;
  assign T_1143 = full == 1'h0;
  assign T_1255 = T_1010 - T_1012;
  assign ptr_diff = T_1255[0:0];
  assign T_1256 = maybe_full & ptr_match;
  assign T_1257 = {T_1256,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_header_src[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_header_dst[initvar] = GEN_1[1:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_addr_beat[initvar] = GEN_2[2:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_client_xact_id[initvar] = GEN_3[0:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_manager_xact_id[initvar] = GEN_4[1:0];
  `endif
  GEN_5 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_is_builtin_type[initvar] = GEN_5[0:0];
  `endif
  GEN_6 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_g_type[initvar] = GEN_6[3:0];
  `endif
  GEN_7 = {2{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_data[initvar] = GEN_7[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_8 = {1{$random}};
  T_1010 = GEN_8[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_9 = {1{$random}};
  T_1012 = GEN_9[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_10 = {1{$random}};
  maybe_full = GEN_10[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_header_src_T_1018_en & ram_header_src_T_1018_mask) begin
      ram_header_src[ram_header_src_T_1018_addr] <= ram_header_src_T_1018_data;
    end
    if(ram_header_dst_T_1018_en & ram_header_dst_T_1018_mask) begin
      ram_header_dst[ram_header_dst_T_1018_addr] <= ram_header_dst_T_1018_data;
    end
    if(ram_payload_addr_beat_T_1018_en & ram_payload_addr_beat_T_1018_mask) begin
      ram_payload_addr_beat[ram_payload_addr_beat_T_1018_addr] <= ram_payload_addr_beat_T_1018_data;
    end
    if(ram_payload_client_xact_id_T_1018_en & ram_payload_client_xact_id_T_1018_mask) begin
      ram_payload_client_xact_id[ram_payload_client_xact_id_T_1018_addr] <= ram_payload_client_xact_id_T_1018_data;
    end
    if(ram_payload_manager_xact_id_T_1018_en & ram_payload_manager_xact_id_T_1018_mask) begin
      ram_payload_manager_xact_id[ram_payload_manager_xact_id_T_1018_addr] <= ram_payload_manager_xact_id_T_1018_data;
    end
    if(ram_payload_is_builtin_type_T_1018_en & ram_payload_is_builtin_type_T_1018_mask) begin
      ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1018_addr] <= ram_payload_is_builtin_type_T_1018_data;
    end
    if(ram_payload_g_type_T_1018_en & ram_payload_g_type_T_1018_mask) begin
      ram_payload_g_type[ram_payload_g_type_T_1018_addr] <= ram_payload_g_type_T_1018_data;
    end
    if(ram_payload_data_T_1018_en & ram_payload_data_T_1018_mask) begin
      ram_payload_data[ram_payload_data_T_1018_addr] <= ram_payload_data_T_1018_data;
    end
    if(reset) begin
      T_1010 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_1010 <= T_1133;
      end
    end
    if(reset) begin
      T_1012 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_1012 <= T_1138;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_1139) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module TileLinkEnqueuer(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [1:0] io_client_acquire_bits_header_src,
  input  [1:0] io_client_acquire_bits_header_dst,
  input  [25:0] io_client_acquire_bits_payload_addr_block,
  input   io_client_acquire_bits_payload_client_xact_id,
  input  [2:0] io_client_acquire_bits_payload_addr_beat,
  input   io_client_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_client_acquire_bits_payload_a_type,
  input  [11:0] io_client_acquire_bits_payload_union,
  input  [63:0] io_client_acquire_bits_payload_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [1:0] io_client_grant_bits_header_src,
  output [1:0] io_client_grant_bits_header_dst,
  output [2:0] io_client_grant_bits_payload_addr_beat,
  output  io_client_grant_bits_payload_client_xact_id,
  output [1:0] io_client_grant_bits_payload_manager_xact_id,
  output  io_client_grant_bits_payload_is_builtin_type,
  output [3:0] io_client_grant_bits_payload_g_type,
  output [63:0] io_client_grant_bits_payload_data,
  output  io_client_finish_ready,
  input   io_client_finish_valid,
  input  [1:0] io_client_finish_bits_header_src,
  input  [1:0] io_client_finish_bits_header_dst,
  input  [1:0] io_client_finish_bits_payload_manager_xact_id,
  input   io_client_probe_ready,
  output  io_client_probe_valid,
  output [1:0] io_client_probe_bits_header_src,
  output [1:0] io_client_probe_bits_header_dst,
  output [25:0] io_client_probe_bits_payload_addr_block,
  output [1:0] io_client_probe_bits_payload_p_type,
  output  io_client_release_ready,
  input   io_client_release_valid,
  input  [1:0] io_client_release_bits_header_src,
  input  [1:0] io_client_release_bits_header_dst,
  input  [2:0] io_client_release_bits_payload_addr_beat,
  input  [25:0] io_client_release_bits_payload_addr_block,
  input   io_client_release_bits_payload_client_xact_id,
  input   io_client_release_bits_payload_voluntary,
  input  [2:0] io_client_release_bits_payload_r_type,
  input  [63:0] io_client_release_bits_payload_data,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [1:0] io_manager_acquire_bits_header_src,
  output [1:0] io_manager_acquire_bits_header_dst,
  output [25:0] io_manager_acquire_bits_payload_addr_block,
  output  io_manager_acquire_bits_payload_client_xact_id,
  output [2:0] io_manager_acquire_bits_payload_addr_beat,
  output  io_manager_acquire_bits_payload_is_builtin_type,
  output [2:0] io_manager_acquire_bits_payload_a_type,
  output [11:0] io_manager_acquire_bits_payload_union,
  output [63:0] io_manager_acquire_bits_payload_data,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [1:0] io_manager_grant_bits_header_src,
  input  [1:0] io_manager_grant_bits_header_dst,
  input  [2:0] io_manager_grant_bits_payload_addr_beat,
  input   io_manager_grant_bits_payload_client_xact_id,
  input  [1:0] io_manager_grant_bits_payload_manager_xact_id,
  input   io_manager_grant_bits_payload_is_builtin_type,
  input  [3:0] io_manager_grant_bits_payload_g_type,
  input  [63:0] io_manager_grant_bits_payload_data,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [1:0] io_manager_finish_bits_header_src,
  output [1:0] io_manager_finish_bits_header_dst,
  output [1:0] io_manager_finish_bits_payload_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [1:0] io_manager_probe_bits_header_src,
  input  [1:0] io_manager_probe_bits_header_dst,
  input  [25:0] io_manager_probe_bits_payload_addr_block,
  input  [1:0] io_manager_probe_bits_payload_p_type,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [1:0] io_manager_release_bits_header_src,
  output [1:0] io_manager_release_bits_header_dst,
  output [2:0] io_manager_release_bits_payload_addr_beat,
  output [25:0] io_manager_release_bits_payload_addr_block,
  output  io_manager_release_bits_payload_client_xact_id,
  output  io_manager_release_bits_payload_voluntary,
  output [2:0] io_manager_release_bits_payload_r_type,
  output [63:0] io_manager_release_bits_payload_data
);
  wire  Queue_4_clk;
  wire  Queue_4_reset;
  wire  Queue_4_io_enq_ready;
  wire  Queue_4_io_enq_valid;
  wire [1:0] Queue_4_io_enq_bits_header_src;
  wire [1:0] Queue_4_io_enq_bits_header_dst;
  wire [25:0] Queue_4_io_enq_bits_payload_addr_block;
  wire  Queue_4_io_enq_bits_payload_client_xact_id;
  wire [2:0] Queue_4_io_enq_bits_payload_addr_beat;
  wire  Queue_4_io_enq_bits_payload_is_builtin_type;
  wire [2:0] Queue_4_io_enq_bits_payload_a_type;
  wire [11:0] Queue_4_io_enq_bits_payload_union;
  wire [63:0] Queue_4_io_enq_bits_payload_data;
  wire  Queue_4_io_deq_ready;
  wire  Queue_4_io_deq_valid;
  wire [1:0] Queue_4_io_deq_bits_header_src;
  wire [1:0] Queue_4_io_deq_bits_header_dst;
  wire [25:0] Queue_4_io_deq_bits_payload_addr_block;
  wire  Queue_4_io_deq_bits_payload_client_xact_id;
  wire [2:0] Queue_4_io_deq_bits_payload_addr_beat;
  wire  Queue_4_io_deq_bits_payload_is_builtin_type;
  wire [2:0] Queue_4_io_deq_bits_payload_a_type;
  wire [11:0] Queue_4_io_deq_bits_payload_union;
  wire [63:0] Queue_4_io_deq_bits_payload_data;
  wire  Queue_4_io_count;
  wire  Queue_1_1_clk;
  wire  Queue_1_1_reset;
  wire  Queue_1_1_io_enq_ready;
  wire  Queue_1_1_io_enq_valid;
  wire [1:0] Queue_1_1_io_enq_bits_header_src;
  wire [1:0] Queue_1_1_io_enq_bits_header_dst;
  wire [25:0] Queue_1_1_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_1_1_io_enq_bits_payload_p_type;
  wire  Queue_1_1_io_deq_ready;
  wire  Queue_1_1_io_deq_valid;
  wire [1:0] Queue_1_1_io_deq_bits_header_src;
  wire [1:0] Queue_1_1_io_deq_bits_header_dst;
  wire [25:0] Queue_1_1_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_1_1_io_deq_bits_payload_p_type;
  wire  Queue_1_1_io_count;
  wire  Queue_2_1_clk;
  wire  Queue_2_1_reset;
  wire  Queue_2_1_io_enq_ready;
  wire  Queue_2_1_io_enq_valid;
  wire [1:0] Queue_2_1_io_enq_bits_header_src;
  wire [1:0] Queue_2_1_io_enq_bits_header_dst;
  wire [2:0] Queue_2_1_io_enq_bits_payload_addr_beat;
  wire [25:0] Queue_2_1_io_enq_bits_payload_addr_block;
  wire  Queue_2_1_io_enq_bits_payload_client_xact_id;
  wire  Queue_2_1_io_enq_bits_payload_voluntary;
  wire [2:0] Queue_2_1_io_enq_bits_payload_r_type;
  wire [63:0] Queue_2_1_io_enq_bits_payload_data;
  wire  Queue_2_1_io_deq_ready;
  wire  Queue_2_1_io_deq_valid;
  wire [1:0] Queue_2_1_io_deq_bits_header_src;
  wire [1:0] Queue_2_1_io_deq_bits_header_dst;
  wire [2:0] Queue_2_1_io_deq_bits_payload_addr_beat;
  wire [25:0] Queue_2_1_io_deq_bits_payload_addr_block;
  wire  Queue_2_1_io_deq_bits_payload_client_xact_id;
  wire  Queue_2_1_io_deq_bits_payload_voluntary;
  wire [2:0] Queue_2_1_io_deq_bits_payload_r_type;
  wire [63:0] Queue_2_1_io_deq_bits_payload_data;
  wire [1:0] Queue_2_1_io_count;
  wire  Queue_3_1_clk;
  wire  Queue_3_1_reset;
  wire  Queue_3_1_io_enq_ready;
  wire  Queue_3_1_io_enq_valid;
  wire [1:0] Queue_3_1_io_enq_bits_header_src;
  wire [1:0] Queue_3_1_io_enq_bits_header_dst;
  wire [2:0] Queue_3_1_io_enq_bits_payload_addr_beat;
  wire  Queue_3_1_io_enq_bits_payload_client_xact_id;
  wire [1:0] Queue_3_1_io_enq_bits_payload_manager_xact_id;
  wire  Queue_3_1_io_enq_bits_payload_is_builtin_type;
  wire [3:0] Queue_3_1_io_enq_bits_payload_g_type;
  wire [63:0] Queue_3_1_io_enq_bits_payload_data;
  wire  Queue_3_1_io_deq_ready;
  wire  Queue_3_1_io_deq_valid;
  wire [1:0] Queue_3_1_io_deq_bits_header_src;
  wire [1:0] Queue_3_1_io_deq_bits_header_dst;
  wire [2:0] Queue_3_1_io_deq_bits_payload_addr_beat;
  wire  Queue_3_1_io_deq_bits_payload_client_xact_id;
  wire [1:0] Queue_3_1_io_deq_bits_payload_manager_xact_id;
  wire  Queue_3_1_io_deq_bits_payload_is_builtin_type;
  wire [3:0] Queue_3_1_io_deq_bits_payload_g_type;
  wire [63:0] Queue_3_1_io_deq_bits_payload_data;
  wire [1:0] Queue_3_1_io_count;
  Queue Queue_4 (
    .clk(Queue_4_clk),
    .reset(Queue_4_reset),
    .io_enq_ready(Queue_4_io_enq_ready),
    .io_enq_valid(Queue_4_io_enq_valid),
    .io_enq_bits_header_src(Queue_4_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_4_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_4_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_4_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_addr_beat(Queue_4_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_is_builtin_type(Queue_4_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_a_type(Queue_4_io_enq_bits_payload_a_type),
    .io_enq_bits_payload_union(Queue_4_io_enq_bits_payload_union),
    .io_enq_bits_payload_data(Queue_4_io_enq_bits_payload_data),
    .io_deq_ready(Queue_4_io_deq_ready),
    .io_deq_valid(Queue_4_io_deq_valid),
    .io_deq_bits_header_src(Queue_4_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_4_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_4_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_4_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_addr_beat(Queue_4_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_is_builtin_type(Queue_4_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_a_type(Queue_4_io_deq_bits_payload_a_type),
    .io_deq_bits_payload_union(Queue_4_io_deq_bits_payload_union),
    .io_deq_bits_payload_data(Queue_4_io_deq_bits_payload_data),
    .io_count(Queue_4_io_count)
  );
  Queue_1 Queue_1_1 (
    .clk(Queue_1_1_clk),
    .reset(Queue_1_1_reset),
    .io_enq_ready(Queue_1_1_io_enq_ready),
    .io_enq_valid(Queue_1_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_1_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_1_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_1_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_p_type(Queue_1_1_io_enq_bits_payload_p_type),
    .io_deq_ready(Queue_1_1_io_deq_ready),
    .io_deq_valid(Queue_1_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_1_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_1_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_1_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_p_type(Queue_1_1_io_deq_bits_payload_p_type),
    .io_count(Queue_1_1_io_count)
  );
  Queue_2 Queue_2_1 (
    .clk(Queue_2_1_clk),
    .reset(Queue_2_1_reset),
    .io_enq_ready(Queue_2_1_io_enq_ready),
    .io_enq_valid(Queue_2_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_2_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_2_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_2_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_addr_block(Queue_2_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_2_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_voluntary(Queue_2_1_io_enq_bits_payload_voluntary),
    .io_enq_bits_payload_r_type(Queue_2_1_io_enq_bits_payload_r_type),
    .io_enq_bits_payload_data(Queue_2_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_2_1_io_deq_ready),
    .io_deq_valid(Queue_2_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_2_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_2_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_2_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_addr_block(Queue_2_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_2_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_voluntary(Queue_2_1_io_deq_bits_payload_voluntary),
    .io_deq_bits_payload_r_type(Queue_2_1_io_deq_bits_payload_r_type),
    .io_deq_bits_payload_data(Queue_2_1_io_deq_bits_payload_data),
    .io_count(Queue_2_1_io_count)
  );
  Queue_3 Queue_3_1 (
    .clk(Queue_3_1_clk),
    .reset(Queue_3_1_reset),
    .io_enq_ready(Queue_3_1_io_enq_ready),
    .io_enq_valid(Queue_3_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_3_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_3_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_3_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_client_xact_id(Queue_3_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_manager_xact_id(Queue_3_1_io_enq_bits_payload_manager_xact_id),
    .io_enq_bits_payload_is_builtin_type(Queue_3_1_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_g_type(Queue_3_1_io_enq_bits_payload_g_type),
    .io_enq_bits_payload_data(Queue_3_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_3_1_io_deq_ready),
    .io_deq_valid(Queue_3_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_3_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_3_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_3_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_client_xact_id(Queue_3_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_manager_xact_id(Queue_3_1_io_deq_bits_payload_manager_xact_id),
    .io_deq_bits_payload_is_builtin_type(Queue_3_1_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_g_type(Queue_3_1_io_deq_bits_payload_g_type),
    .io_deq_bits_payload_data(Queue_3_1_io_deq_bits_payload_data),
    .io_count(Queue_3_1_io_count)
  );
  assign io_client_acquire_ready = Queue_4_io_enq_ready;
  assign io_client_grant_valid = Queue_3_1_io_deq_valid;
  assign io_client_grant_bits_header_src = Queue_3_1_io_deq_bits_header_src;
  assign io_client_grant_bits_header_dst = Queue_3_1_io_deq_bits_header_dst;
  assign io_client_grant_bits_payload_addr_beat = Queue_3_1_io_deq_bits_payload_addr_beat;
  assign io_client_grant_bits_payload_client_xact_id = Queue_3_1_io_deq_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_manager_xact_id = Queue_3_1_io_deq_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_is_builtin_type = Queue_3_1_io_deq_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_g_type = Queue_3_1_io_deq_bits_payload_g_type;
  assign io_client_grant_bits_payload_data = Queue_3_1_io_deq_bits_payload_data;
  assign io_client_finish_ready = io_manager_finish_ready;
  assign io_client_probe_valid = Queue_1_1_io_deq_valid;
  assign io_client_probe_bits_header_src = Queue_1_1_io_deq_bits_header_src;
  assign io_client_probe_bits_header_dst = Queue_1_1_io_deq_bits_header_dst;
  assign io_client_probe_bits_payload_addr_block = Queue_1_1_io_deq_bits_payload_addr_block;
  assign io_client_probe_bits_payload_p_type = Queue_1_1_io_deq_bits_payload_p_type;
  assign io_client_release_ready = Queue_2_1_io_enq_ready;
  assign io_manager_acquire_valid = Queue_4_io_deq_valid;
  assign io_manager_acquire_bits_header_src = Queue_4_io_deq_bits_header_src;
  assign io_manager_acquire_bits_header_dst = Queue_4_io_deq_bits_header_dst;
  assign io_manager_acquire_bits_payload_addr_block = Queue_4_io_deq_bits_payload_addr_block;
  assign io_manager_acquire_bits_payload_client_xact_id = Queue_4_io_deq_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_beat = Queue_4_io_deq_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_is_builtin_type = Queue_4_io_deq_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_a_type = Queue_4_io_deq_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_union = Queue_4_io_deq_bits_payload_union;
  assign io_manager_acquire_bits_payload_data = Queue_4_io_deq_bits_payload_data;
  assign io_manager_grant_ready = Queue_3_1_io_enq_ready;
  assign io_manager_finish_valid = io_client_finish_valid;
  assign io_manager_finish_bits_header_src = io_client_finish_bits_header_src;
  assign io_manager_finish_bits_header_dst = io_client_finish_bits_header_dst;
  assign io_manager_finish_bits_payload_manager_xact_id = io_client_finish_bits_payload_manager_xact_id;
  assign io_manager_probe_ready = Queue_1_1_io_enq_ready;
  assign io_manager_release_valid = Queue_2_1_io_deq_valid;
  assign io_manager_release_bits_header_src = Queue_2_1_io_deq_bits_header_src;
  assign io_manager_release_bits_header_dst = Queue_2_1_io_deq_bits_header_dst;
  assign io_manager_release_bits_payload_addr_beat = Queue_2_1_io_deq_bits_payload_addr_beat;
  assign io_manager_release_bits_payload_addr_block = Queue_2_1_io_deq_bits_payload_addr_block;
  assign io_manager_release_bits_payload_client_xact_id = Queue_2_1_io_deq_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_voluntary = Queue_2_1_io_deq_bits_payload_voluntary;
  assign io_manager_release_bits_payload_r_type = Queue_2_1_io_deq_bits_payload_r_type;
  assign io_manager_release_bits_payload_data = Queue_2_1_io_deq_bits_payload_data;
  assign Queue_4_clk = clk;
  assign Queue_4_reset = reset;
  assign Queue_4_io_enq_valid = io_client_acquire_valid;
  assign Queue_4_io_enq_bits_header_src = io_client_acquire_bits_header_src;
  assign Queue_4_io_enq_bits_header_dst = io_client_acquire_bits_header_dst;
  assign Queue_4_io_enq_bits_payload_addr_block = io_client_acquire_bits_payload_addr_block;
  assign Queue_4_io_enq_bits_payload_client_xact_id = io_client_acquire_bits_payload_client_xact_id;
  assign Queue_4_io_enq_bits_payload_addr_beat = io_client_acquire_bits_payload_addr_beat;
  assign Queue_4_io_enq_bits_payload_is_builtin_type = io_client_acquire_bits_payload_is_builtin_type;
  assign Queue_4_io_enq_bits_payload_a_type = io_client_acquire_bits_payload_a_type;
  assign Queue_4_io_enq_bits_payload_union = io_client_acquire_bits_payload_union;
  assign Queue_4_io_enq_bits_payload_data = io_client_acquire_bits_payload_data;
  assign Queue_4_io_deq_ready = io_manager_acquire_ready;
  assign Queue_1_1_clk = clk;
  assign Queue_1_1_reset = reset;
  assign Queue_1_1_io_enq_valid = io_manager_probe_valid;
  assign Queue_1_1_io_enq_bits_header_src = io_manager_probe_bits_header_src;
  assign Queue_1_1_io_enq_bits_header_dst = io_manager_probe_bits_header_dst;
  assign Queue_1_1_io_enq_bits_payload_addr_block = io_manager_probe_bits_payload_addr_block;
  assign Queue_1_1_io_enq_bits_payload_p_type = io_manager_probe_bits_payload_p_type;
  assign Queue_1_1_io_deq_ready = io_client_probe_ready;
  assign Queue_2_1_clk = clk;
  assign Queue_2_1_reset = reset;
  assign Queue_2_1_io_enq_valid = io_client_release_valid;
  assign Queue_2_1_io_enq_bits_header_src = io_client_release_bits_header_src;
  assign Queue_2_1_io_enq_bits_header_dst = io_client_release_bits_header_dst;
  assign Queue_2_1_io_enq_bits_payload_addr_beat = io_client_release_bits_payload_addr_beat;
  assign Queue_2_1_io_enq_bits_payload_addr_block = io_client_release_bits_payload_addr_block;
  assign Queue_2_1_io_enq_bits_payload_client_xact_id = io_client_release_bits_payload_client_xact_id;
  assign Queue_2_1_io_enq_bits_payload_voluntary = io_client_release_bits_payload_voluntary;
  assign Queue_2_1_io_enq_bits_payload_r_type = io_client_release_bits_payload_r_type;
  assign Queue_2_1_io_enq_bits_payload_data = io_client_release_bits_payload_data;
  assign Queue_2_1_io_deq_ready = io_manager_release_ready;
  assign Queue_3_1_clk = clk;
  assign Queue_3_1_reset = reset;
  assign Queue_3_1_io_enq_valid = io_manager_grant_valid;
  assign Queue_3_1_io_enq_bits_header_src = io_manager_grant_bits_header_src;
  assign Queue_3_1_io_enq_bits_header_dst = io_manager_grant_bits_header_dst;
  assign Queue_3_1_io_enq_bits_payload_addr_beat = io_manager_grant_bits_payload_addr_beat;
  assign Queue_3_1_io_enq_bits_payload_client_xact_id = io_manager_grant_bits_payload_client_xact_id;
  assign Queue_3_1_io_enq_bits_payload_manager_xact_id = io_manager_grant_bits_payload_manager_xact_id;
  assign Queue_3_1_io_enq_bits_payload_is_builtin_type = io_manager_grant_bits_payload_is_builtin_type;
  assign Queue_3_1_io_enq_bits_payload_g_type = io_manager_grant_bits_payload_g_type;
  assign Queue_3_1_io_enq_bits_payload_data = io_manager_grant_bits_payload_data;
  assign Queue_3_1_io_deq_ready = io_client_grant_ready;
endmodule
module ClientTileLinkNetworkPort(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [25:0] io_client_acquire_bits_addr_block,
  input   io_client_acquire_bits_client_xact_id,
  input  [2:0] io_client_acquire_bits_addr_beat,
  input   io_client_acquire_bits_is_builtin_type,
  input  [2:0] io_client_acquire_bits_a_type,
  input  [11:0] io_client_acquire_bits_union,
  input  [63:0] io_client_acquire_bits_data,
  input   io_client_probe_ready,
  output  io_client_probe_valid,
  output [25:0] io_client_probe_bits_addr_block,
  output [1:0] io_client_probe_bits_p_type,
  output  io_client_release_ready,
  input   io_client_release_valid,
  input  [2:0] io_client_release_bits_addr_beat,
  input  [25:0] io_client_release_bits_addr_block,
  input   io_client_release_bits_client_xact_id,
  input   io_client_release_bits_voluntary,
  input  [2:0] io_client_release_bits_r_type,
  input  [63:0] io_client_release_bits_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [2:0] io_client_grant_bits_addr_beat,
  output  io_client_grant_bits_client_xact_id,
  output [1:0] io_client_grant_bits_manager_xact_id,
  output  io_client_grant_bits_is_builtin_type,
  output [3:0] io_client_grant_bits_g_type,
  output [63:0] io_client_grant_bits_data,
  output  io_client_grant_bits_manager_id,
  output  io_client_finish_ready,
  input   io_client_finish_valid,
  input  [1:0] io_client_finish_bits_manager_xact_id,
  input   io_client_finish_bits_manager_id,
  input   io_network_acquire_ready,
  output  io_network_acquire_valid,
  output [1:0] io_network_acquire_bits_header_src,
  output [1:0] io_network_acquire_bits_header_dst,
  output [25:0] io_network_acquire_bits_payload_addr_block,
  output  io_network_acquire_bits_payload_client_xact_id,
  output [2:0] io_network_acquire_bits_payload_addr_beat,
  output  io_network_acquire_bits_payload_is_builtin_type,
  output [2:0] io_network_acquire_bits_payload_a_type,
  output [11:0] io_network_acquire_bits_payload_union,
  output [63:0] io_network_acquire_bits_payload_data,
  output  io_network_grant_ready,
  input   io_network_grant_valid,
  input  [1:0] io_network_grant_bits_header_src,
  input  [1:0] io_network_grant_bits_header_dst,
  input  [2:0] io_network_grant_bits_payload_addr_beat,
  input   io_network_grant_bits_payload_client_xact_id,
  input  [1:0] io_network_grant_bits_payload_manager_xact_id,
  input   io_network_grant_bits_payload_is_builtin_type,
  input  [3:0] io_network_grant_bits_payload_g_type,
  input  [63:0] io_network_grant_bits_payload_data,
  input   io_network_finish_ready,
  output  io_network_finish_valid,
  output [1:0] io_network_finish_bits_header_src,
  output [1:0] io_network_finish_bits_header_dst,
  output [1:0] io_network_finish_bits_payload_manager_xact_id,
  output  io_network_probe_ready,
  input   io_network_probe_valid,
  input  [1:0] io_network_probe_bits_header_src,
  input  [1:0] io_network_probe_bits_header_dst,
  input  [25:0] io_network_probe_bits_payload_addr_block,
  input  [1:0] io_network_probe_bits_payload_p_type,
  input   io_network_release_ready,
  output  io_network_release_valid,
  output [1:0] io_network_release_bits_header_src,
  output [1:0] io_network_release_bits_header_dst,
  output [2:0] io_network_release_bits_payload_addr_beat,
  output [25:0] io_network_release_bits_payload_addr_block,
  output  io_network_release_bits_payload_client_xact_id,
  output  io_network_release_bits_payload_voluntary,
  output [2:0] io_network_release_bits_payload_r_type,
  output [63:0] io_network_release_bits_payload_data
);
  wire  acq_with_header_ready;
  wire  acq_with_header_valid;
  wire [1:0] acq_with_header_bits_header_src;
  wire [1:0] acq_with_header_bits_header_dst;
  wire [25:0] acq_with_header_bits_payload_addr_block;
  wire  acq_with_header_bits_payload_client_xact_id;
  wire [2:0] acq_with_header_bits_payload_addr_beat;
  wire  acq_with_header_bits_payload_is_builtin_type;
  wire [2:0] acq_with_header_bits_payload_a_type;
  wire [11:0] acq_with_header_bits_payload_union;
  wire [63:0] acq_with_header_bits_payload_data;
  wire [31:0] GEN_0;
  wire [31:0] T_3894;
  wire  T_3896;
  wire  T_3898;
  wire  T_3899;
  wire  T_3902;
  wire  rel_with_header_ready;
  wire  rel_with_header_valid;
  wire [1:0] rel_with_header_bits_header_src;
  wire [1:0] rel_with_header_bits_header_dst;
  wire [2:0] rel_with_header_bits_payload_addr_beat;
  wire [25:0] rel_with_header_bits_payload_addr_block;
  wire  rel_with_header_bits_payload_client_xact_id;
  wire  rel_with_header_bits_payload_voluntary;
  wire [2:0] rel_with_header_bits_payload_r_type;
  wire [63:0] rel_with_header_bits_payload_data;
  wire [31:0] GEN_1;
  wire [31:0] T_4464;
  wire  T_4466;
  wire  T_4468;
  wire  T_4469;
  wire  T_4472;
  wire  fin_with_header_ready;
  wire  fin_with_header_valid;
  wire [1:0] fin_with_header_bits_header_src;
  wire [1:0] fin_with_header_bits_header_dst;
  wire [1:0] fin_with_header_bits_payload_manager_xact_id;
  wire  fin_with_header_bits_payload_manager_id;
  wire  prb_without_header_ready;
  wire  prb_without_header_valid;
  wire [25:0] prb_without_header_bits_addr_block;
  wire [1:0] prb_without_header_bits_p_type;
  wire  gnt_without_header_ready;
  wire  gnt_without_header_valid;
  wire [2:0] gnt_without_header_bits_addr_beat;
  wire  gnt_without_header_bits_client_xact_id;
  wire [1:0] gnt_without_header_bits_manager_xact_id;
  wire  gnt_without_header_bits_is_builtin_type;
  wire [3:0] gnt_without_header_bits_g_type;
  wire [63:0] gnt_without_header_bits_data;
  assign io_client_acquire_ready = acq_with_header_ready;
  assign io_client_probe_valid = prb_without_header_valid;
  assign io_client_probe_bits_addr_block = prb_without_header_bits_addr_block;
  assign io_client_probe_bits_p_type = prb_without_header_bits_p_type;
  assign io_client_release_ready = rel_with_header_ready;
  assign io_client_grant_valid = gnt_without_header_valid;
  assign io_client_grant_bits_addr_beat = gnt_without_header_bits_addr_beat;
  assign io_client_grant_bits_client_xact_id = gnt_without_header_bits_client_xact_id;
  assign io_client_grant_bits_manager_xact_id = gnt_without_header_bits_manager_xact_id;
  assign io_client_grant_bits_is_builtin_type = gnt_without_header_bits_is_builtin_type;
  assign io_client_grant_bits_g_type = gnt_without_header_bits_g_type;
  assign io_client_grant_bits_data = gnt_without_header_bits_data;
  assign io_client_grant_bits_manager_id = io_network_grant_bits_header_src[0];
  assign io_client_finish_ready = fin_with_header_ready;
  assign io_network_acquire_valid = acq_with_header_valid;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign io_network_grant_ready = gnt_without_header_ready;
  assign io_network_finish_valid = fin_with_header_valid;
  assign io_network_finish_bits_header_src = fin_with_header_bits_header_src;
  assign io_network_finish_bits_header_dst = fin_with_header_bits_header_dst;
  assign io_network_finish_bits_payload_manager_xact_id = fin_with_header_bits_payload_manager_xact_id;
  assign io_network_probe_ready = prb_without_header_ready;
  assign io_network_release_valid = rel_with_header_valid;
  assign io_network_release_bits_header_src = rel_with_header_bits_header_src;
  assign io_network_release_bits_header_dst = rel_with_header_bits_header_dst;
  assign io_network_release_bits_payload_addr_beat = rel_with_header_bits_payload_addr_beat;
  assign io_network_release_bits_payload_addr_block = rel_with_header_bits_payload_addr_block;
  assign io_network_release_bits_payload_client_xact_id = rel_with_header_bits_payload_client_xact_id;
  assign io_network_release_bits_payload_voluntary = rel_with_header_bits_payload_voluntary;
  assign io_network_release_bits_payload_r_type = rel_with_header_bits_payload_r_type;
  assign io_network_release_bits_payload_data = rel_with_header_bits_payload_data;
  assign acq_with_header_ready = io_network_acquire_ready;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign acq_with_header_bits_header_src = 2'h0;
  assign acq_with_header_bits_header_dst = {{1'd0}, T_3902};
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign GEN_0 = {{6'd0}, io_client_acquire_bits_addr_block};
  assign T_3894 = GEN_0 << 6;
  assign T_3896 = 32'h80000000 <= T_3894;
  assign T_3898 = T_3894 < 32'h90000000;
  assign T_3899 = T_3896 & T_3898;
  assign T_3902 = T_3899 ? 1'h0 : 1'h1;
  assign rel_with_header_ready = io_network_release_ready;
  assign rel_with_header_valid = io_client_release_valid;
  assign rel_with_header_bits_header_src = 2'h0;
  assign rel_with_header_bits_header_dst = {{1'd0}, T_4472};
  assign rel_with_header_bits_payload_addr_beat = io_client_release_bits_addr_beat;
  assign rel_with_header_bits_payload_addr_block = io_client_release_bits_addr_block;
  assign rel_with_header_bits_payload_client_xact_id = io_client_release_bits_client_xact_id;
  assign rel_with_header_bits_payload_voluntary = io_client_release_bits_voluntary;
  assign rel_with_header_bits_payload_r_type = io_client_release_bits_r_type;
  assign rel_with_header_bits_payload_data = io_client_release_bits_data;
  assign GEN_1 = {{6'd0}, io_client_release_bits_addr_block};
  assign T_4464 = GEN_1 << 6;
  assign T_4466 = 32'h80000000 <= T_4464;
  assign T_4468 = T_4464 < 32'h90000000;
  assign T_4469 = T_4466 & T_4468;
  assign T_4472 = T_4469 ? 1'h0 : 1'h1;
  assign fin_with_header_ready = io_network_finish_ready;
  assign fin_with_header_valid = io_client_finish_valid;
  assign fin_with_header_bits_header_src = 2'h0;
  assign fin_with_header_bits_header_dst = {{1'd0}, io_client_finish_bits_manager_id};
  assign fin_with_header_bits_payload_manager_xact_id = io_client_finish_bits_manager_xact_id;
  assign fin_with_header_bits_payload_manager_id = io_client_finish_bits_manager_id;
  assign prb_without_header_ready = io_client_probe_ready;
  assign prb_without_header_valid = io_network_probe_valid;
  assign prb_without_header_bits_addr_block = io_network_probe_bits_payload_addr_block;
  assign prb_without_header_bits_p_type = io_network_probe_bits_payload_p_type;
  assign gnt_without_header_ready = io_client_grant_ready;
  assign gnt_without_header_valid = io_network_grant_valid;
  assign gnt_without_header_bits_addr_beat = io_network_grant_bits_payload_addr_beat;
  assign gnt_without_header_bits_client_xact_id = io_network_grant_bits_payload_client_xact_id;
  assign gnt_without_header_bits_manager_xact_id = io_network_grant_bits_payload_manager_xact_id;
  assign gnt_without_header_bits_is_builtin_type = io_network_grant_bits_payload_is_builtin_type;
  assign gnt_without_header_bits_g_type = io_network_grant_bits_payload_g_type;
  assign gnt_without_header_bits_data = io_network_grant_bits_payload_data;
endmodule
module TileLinkEnqueuer_1(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [1:0] io_client_acquire_bits_header_src,
  input  [1:0] io_client_acquire_bits_header_dst,
  input  [25:0] io_client_acquire_bits_payload_addr_block,
  input   io_client_acquire_bits_payload_client_xact_id,
  input  [2:0] io_client_acquire_bits_payload_addr_beat,
  input   io_client_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_client_acquire_bits_payload_a_type,
  input  [11:0] io_client_acquire_bits_payload_union,
  input  [63:0] io_client_acquire_bits_payload_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [1:0] io_client_grant_bits_header_src,
  output [1:0] io_client_grant_bits_header_dst,
  output [2:0] io_client_grant_bits_payload_addr_beat,
  output  io_client_grant_bits_payload_client_xact_id,
  output [1:0] io_client_grant_bits_payload_manager_xact_id,
  output  io_client_grant_bits_payload_is_builtin_type,
  output [3:0] io_client_grant_bits_payload_g_type,
  output [63:0] io_client_grant_bits_payload_data,
  output  io_client_finish_ready,
  input   io_client_finish_valid,
  input  [1:0] io_client_finish_bits_header_src,
  input  [1:0] io_client_finish_bits_header_dst,
  input  [1:0] io_client_finish_bits_payload_manager_xact_id,
  input   io_client_probe_ready,
  output  io_client_probe_valid,
  output [1:0] io_client_probe_bits_header_src,
  output [1:0] io_client_probe_bits_header_dst,
  output [25:0] io_client_probe_bits_payload_addr_block,
  output [1:0] io_client_probe_bits_payload_p_type,
  output  io_client_release_ready,
  input   io_client_release_valid,
  input  [1:0] io_client_release_bits_header_src,
  input  [1:0] io_client_release_bits_header_dst,
  input  [2:0] io_client_release_bits_payload_addr_beat,
  input  [25:0] io_client_release_bits_payload_addr_block,
  input   io_client_release_bits_payload_client_xact_id,
  input   io_client_release_bits_payload_voluntary,
  input  [2:0] io_client_release_bits_payload_r_type,
  input  [63:0] io_client_release_bits_payload_data,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [1:0] io_manager_acquire_bits_header_src,
  output [1:0] io_manager_acquire_bits_header_dst,
  output [25:0] io_manager_acquire_bits_payload_addr_block,
  output  io_manager_acquire_bits_payload_client_xact_id,
  output [2:0] io_manager_acquire_bits_payload_addr_beat,
  output  io_manager_acquire_bits_payload_is_builtin_type,
  output [2:0] io_manager_acquire_bits_payload_a_type,
  output [11:0] io_manager_acquire_bits_payload_union,
  output [63:0] io_manager_acquire_bits_payload_data,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [1:0] io_manager_grant_bits_header_src,
  input  [1:0] io_manager_grant_bits_header_dst,
  input  [2:0] io_manager_grant_bits_payload_addr_beat,
  input   io_manager_grant_bits_payload_client_xact_id,
  input  [1:0] io_manager_grant_bits_payload_manager_xact_id,
  input   io_manager_grant_bits_payload_is_builtin_type,
  input  [3:0] io_manager_grant_bits_payload_g_type,
  input  [63:0] io_manager_grant_bits_payload_data,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [1:0] io_manager_finish_bits_header_src,
  output [1:0] io_manager_finish_bits_header_dst,
  output [1:0] io_manager_finish_bits_payload_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [1:0] io_manager_probe_bits_header_src,
  input  [1:0] io_manager_probe_bits_header_dst,
  input  [25:0] io_manager_probe_bits_payload_addr_block,
  input  [1:0] io_manager_probe_bits_payload_p_type,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [1:0] io_manager_release_bits_header_src,
  output [1:0] io_manager_release_bits_header_dst,
  output [2:0] io_manager_release_bits_payload_addr_beat,
  output [25:0] io_manager_release_bits_payload_addr_block,
  output  io_manager_release_bits_payload_client_xact_id,
  output  io_manager_release_bits_payload_voluntary,
  output [2:0] io_manager_release_bits_payload_r_type,
  output [63:0] io_manager_release_bits_payload_data
);
  wire  Queue_4_1_clk;
  wire  Queue_4_1_reset;
  wire  Queue_4_1_io_enq_ready;
  wire  Queue_4_1_io_enq_valid;
  wire [1:0] Queue_4_1_io_enq_bits_header_src;
  wire [1:0] Queue_4_1_io_enq_bits_header_dst;
  wire [25:0] Queue_4_1_io_enq_bits_payload_addr_block;
  wire  Queue_4_1_io_enq_bits_payload_client_xact_id;
  wire [2:0] Queue_4_1_io_enq_bits_payload_addr_beat;
  wire  Queue_4_1_io_enq_bits_payload_is_builtin_type;
  wire [2:0] Queue_4_1_io_enq_bits_payload_a_type;
  wire [11:0] Queue_4_1_io_enq_bits_payload_union;
  wire [63:0] Queue_4_1_io_enq_bits_payload_data;
  wire  Queue_4_1_io_deq_ready;
  wire  Queue_4_1_io_deq_valid;
  wire [1:0] Queue_4_1_io_deq_bits_header_src;
  wire [1:0] Queue_4_1_io_deq_bits_header_dst;
  wire [25:0] Queue_4_1_io_deq_bits_payload_addr_block;
  wire  Queue_4_1_io_deq_bits_payload_client_xact_id;
  wire [2:0] Queue_4_1_io_deq_bits_payload_addr_beat;
  wire  Queue_4_1_io_deq_bits_payload_is_builtin_type;
  wire [2:0] Queue_4_1_io_deq_bits_payload_a_type;
  wire [11:0] Queue_4_1_io_deq_bits_payload_union;
  wire [63:0] Queue_4_1_io_deq_bits_payload_data;
  wire  Queue_4_1_io_count;
  wire  Queue_5_1_clk;
  wire  Queue_5_1_reset;
  wire  Queue_5_1_io_enq_ready;
  wire  Queue_5_1_io_enq_valid;
  wire [1:0] Queue_5_1_io_enq_bits_header_src;
  wire [1:0] Queue_5_1_io_enq_bits_header_dst;
  wire [25:0] Queue_5_1_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_5_1_io_enq_bits_payload_p_type;
  wire  Queue_5_1_io_deq_ready;
  wire  Queue_5_1_io_deq_valid;
  wire [1:0] Queue_5_1_io_deq_bits_header_src;
  wire [1:0] Queue_5_1_io_deq_bits_header_dst;
  wire [25:0] Queue_5_1_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_5_1_io_deq_bits_payload_p_type;
  wire  Queue_5_1_io_count;
  wire  Queue_6_1_clk;
  wire  Queue_6_1_reset;
  wire  Queue_6_1_io_enq_ready;
  wire  Queue_6_1_io_enq_valid;
  wire [1:0] Queue_6_1_io_enq_bits_header_src;
  wire [1:0] Queue_6_1_io_enq_bits_header_dst;
  wire [2:0] Queue_6_1_io_enq_bits_payload_addr_beat;
  wire [25:0] Queue_6_1_io_enq_bits_payload_addr_block;
  wire  Queue_6_1_io_enq_bits_payload_client_xact_id;
  wire  Queue_6_1_io_enq_bits_payload_voluntary;
  wire [2:0] Queue_6_1_io_enq_bits_payload_r_type;
  wire [63:0] Queue_6_1_io_enq_bits_payload_data;
  wire  Queue_6_1_io_deq_ready;
  wire  Queue_6_1_io_deq_valid;
  wire [1:0] Queue_6_1_io_deq_bits_header_src;
  wire [1:0] Queue_6_1_io_deq_bits_header_dst;
  wire [2:0] Queue_6_1_io_deq_bits_payload_addr_beat;
  wire [25:0] Queue_6_1_io_deq_bits_payload_addr_block;
  wire  Queue_6_1_io_deq_bits_payload_client_xact_id;
  wire  Queue_6_1_io_deq_bits_payload_voluntary;
  wire [2:0] Queue_6_1_io_deq_bits_payload_r_type;
  wire [63:0] Queue_6_1_io_deq_bits_payload_data;
  wire [1:0] Queue_6_1_io_count;
  wire  Queue_7_1_clk;
  wire  Queue_7_1_reset;
  wire  Queue_7_1_io_enq_ready;
  wire  Queue_7_1_io_enq_valid;
  wire [1:0] Queue_7_1_io_enq_bits_header_src;
  wire [1:0] Queue_7_1_io_enq_bits_header_dst;
  wire [2:0] Queue_7_1_io_enq_bits_payload_addr_beat;
  wire  Queue_7_1_io_enq_bits_payload_client_xact_id;
  wire [1:0] Queue_7_1_io_enq_bits_payload_manager_xact_id;
  wire  Queue_7_1_io_enq_bits_payload_is_builtin_type;
  wire [3:0] Queue_7_1_io_enq_bits_payload_g_type;
  wire [63:0] Queue_7_1_io_enq_bits_payload_data;
  wire  Queue_7_1_io_deq_ready;
  wire  Queue_7_1_io_deq_valid;
  wire [1:0] Queue_7_1_io_deq_bits_header_src;
  wire [1:0] Queue_7_1_io_deq_bits_header_dst;
  wire [2:0] Queue_7_1_io_deq_bits_payload_addr_beat;
  wire  Queue_7_1_io_deq_bits_payload_client_xact_id;
  wire [1:0] Queue_7_1_io_deq_bits_payload_manager_xact_id;
  wire  Queue_7_1_io_deq_bits_payload_is_builtin_type;
  wire [3:0] Queue_7_1_io_deq_bits_payload_g_type;
  wire [63:0] Queue_7_1_io_deq_bits_payload_data;
  wire [1:0] Queue_7_1_io_count;
  Queue Queue_4_1 (
    .clk(Queue_4_1_clk),
    .reset(Queue_4_1_reset),
    .io_enq_ready(Queue_4_1_io_enq_ready),
    .io_enq_valid(Queue_4_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_4_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_4_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_4_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_4_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_addr_beat(Queue_4_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_is_builtin_type(Queue_4_1_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_a_type(Queue_4_1_io_enq_bits_payload_a_type),
    .io_enq_bits_payload_union(Queue_4_1_io_enq_bits_payload_union),
    .io_enq_bits_payload_data(Queue_4_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_4_1_io_deq_ready),
    .io_deq_valid(Queue_4_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_4_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_4_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_4_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_4_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_addr_beat(Queue_4_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_is_builtin_type(Queue_4_1_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_a_type(Queue_4_1_io_deq_bits_payload_a_type),
    .io_deq_bits_payload_union(Queue_4_1_io_deq_bits_payload_union),
    .io_deq_bits_payload_data(Queue_4_1_io_deq_bits_payload_data),
    .io_count(Queue_4_1_io_count)
  );
  Queue_1 Queue_5_1 (
    .clk(Queue_5_1_clk),
    .reset(Queue_5_1_reset),
    .io_enq_ready(Queue_5_1_io_enq_ready),
    .io_enq_valid(Queue_5_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_5_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_5_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_5_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_p_type(Queue_5_1_io_enq_bits_payload_p_type),
    .io_deq_ready(Queue_5_1_io_deq_ready),
    .io_deq_valid(Queue_5_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_5_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_5_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_5_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_p_type(Queue_5_1_io_deq_bits_payload_p_type),
    .io_count(Queue_5_1_io_count)
  );
  Queue_2 Queue_6_1 (
    .clk(Queue_6_1_clk),
    .reset(Queue_6_1_reset),
    .io_enq_ready(Queue_6_1_io_enq_ready),
    .io_enq_valid(Queue_6_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_6_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_6_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_6_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_addr_block(Queue_6_1_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_6_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_voluntary(Queue_6_1_io_enq_bits_payload_voluntary),
    .io_enq_bits_payload_r_type(Queue_6_1_io_enq_bits_payload_r_type),
    .io_enq_bits_payload_data(Queue_6_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_6_1_io_deq_ready),
    .io_deq_valid(Queue_6_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_6_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_6_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_6_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_addr_block(Queue_6_1_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_6_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_voluntary(Queue_6_1_io_deq_bits_payload_voluntary),
    .io_deq_bits_payload_r_type(Queue_6_1_io_deq_bits_payload_r_type),
    .io_deq_bits_payload_data(Queue_6_1_io_deq_bits_payload_data),
    .io_count(Queue_6_1_io_count)
  );
  Queue_3 Queue_7_1 (
    .clk(Queue_7_1_clk),
    .reset(Queue_7_1_reset),
    .io_enq_ready(Queue_7_1_io_enq_ready),
    .io_enq_valid(Queue_7_1_io_enq_valid),
    .io_enq_bits_header_src(Queue_7_1_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_7_1_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_7_1_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_client_xact_id(Queue_7_1_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_manager_xact_id(Queue_7_1_io_enq_bits_payload_manager_xact_id),
    .io_enq_bits_payload_is_builtin_type(Queue_7_1_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_g_type(Queue_7_1_io_enq_bits_payload_g_type),
    .io_enq_bits_payload_data(Queue_7_1_io_enq_bits_payload_data),
    .io_deq_ready(Queue_7_1_io_deq_ready),
    .io_deq_valid(Queue_7_1_io_deq_valid),
    .io_deq_bits_header_src(Queue_7_1_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_7_1_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_7_1_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_client_xact_id(Queue_7_1_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_manager_xact_id(Queue_7_1_io_deq_bits_payload_manager_xact_id),
    .io_deq_bits_payload_is_builtin_type(Queue_7_1_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_g_type(Queue_7_1_io_deq_bits_payload_g_type),
    .io_deq_bits_payload_data(Queue_7_1_io_deq_bits_payload_data),
    .io_count(Queue_7_1_io_count)
  );
  assign io_client_acquire_ready = Queue_4_1_io_enq_ready;
  assign io_client_grant_valid = Queue_7_1_io_deq_valid;
  assign io_client_grant_bits_header_src = Queue_7_1_io_deq_bits_header_src;
  assign io_client_grant_bits_header_dst = Queue_7_1_io_deq_bits_header_dst;
  assign io_client_grant_bits_payload_addr_beat = Queue_7_1_io_deq_bits_payload_addr_beat;
  assign io_client_grant_bits_payload_client_xact_id = Queue_7_1_io_deq_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_manager_xact_id = Queue_7_1_io_deq_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_is_builtin_type = Queue_7_1_io_deq_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_g_type = Queue_7_1_io_deq_bits_payload_g_type;
  assign io_client_grant_bits_payload_data = Queue_7_1_io_deq_bits_payload_data;
  assign io_client_finish_ready = io_manager_finish_ready;
  assign io_client_probe_valid = Queue_5_1_io_deq_valid;
  assign io_client_probe_bits_header_src = Queue_5_1_io_deq_bits_header_src;
  assign io_client_probe_bits_header_dst = Queue_5_1_io_deq_bits_header_dst;
  assign io_client_probe_bits_payload_addr_block = Queue_5_1_io_deq_bits_payload_addr_block;
  assign io_client_probe_bits_payload_p_type = Queue_5_1_io_deq_bits_payload_p_type;
  assign io_client_release_ready = Queue_6_1_io_enq_ready;
  assign io_manager_acquire_valid = Queue_4_1_io_deq_valid;
  assign io_manager_acquire_bits_header_src = Queue_4_1_io_deq_bits_header_src;
  assign io_manager_acquire_bits_header_dst = Queue_4_1_io_deq_bits_header_dst;
  assign io_manager_acquire_bits_payload_addr_block = Queue_4_1_io_deq_bits_payload_addr_block;
  assign io_manager_acquire_bits_payload_client_xact_id = Queue_4_1_io_deq_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_beat = Queue_4_1_io_deq_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_is_builtin_type = Queue_4_1_io_deq_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_a_type = Queue_4_1_io_deq_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_union = Queue_4_1_io_deq_bits_payload_union;
  assign io_manager_acquire_bits_payload_data = Queue_4_1_io_deq_bits_payload_data;
  assign io_manager_grant_ready = Queue_7_1_io_enq_ready;
  assign io_manager_finish_valid = io_client_finish_valid;
  assign io_manager_finish_bits_header_src = io_client_finish_bits_header_src;
  assign io_manager_finish_bits_header_dst = io_client_finish_bits_header_dst;
  assign io_manager_finish_bits_payload_manager_xact_id = io_client_finish_bits_payload_manager_xact_id;
  assign io_manager_probe_ready = Queue_5_1_io_enq_ready;
  assign io_manager_release_valid = Queue_6_1_io_deq_valid;
  assign io_manager_release_bits_header_src = Queue_6_1_io_deq_bits_header_src;
  assign io_manager_release_bits_header_dst = Queue_6_1_io_deq_bits_header_dst;
  assign io_manager_release_bits_payload_addr_beat = Queue_6_1_io_deq_bits_payload_addr_beat;
  assign io_manager_release_bits_payload_addr_block = Queue_6_1_io_deq_bits_payload_addr_block;
  assign io_manager_release_bits_payload_client_xact_id = Queue_6_1_io_deq_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_voluntary = Queue_6_1_io_deq_bits_payload_voluntary;
  assign io_manager_release_bits_payload_r_type = Queue_6_1_io_deq_bits_payload_r_type;
  assign io_manager_release_bits_payload_data = Queue_6_1_io_deq_bits_payload_data;
  assign Queue_4_1_clk = clk;
  assign Queue_4_1_reset = reset;
  assign Queue_4_1_io_enq_valid = io_client_acquire_valid;
  assign Queue_4_1_io_enq_bits_header_src = io_client_acquire_bits_header_src;
  assign Queue_4_1_io_enq_bits_header_dst = io_client_acquire_bits_header_dst;
  assign Queue_4_1_io_enq_bits_payload_addr_block = io_client_acquire_bits_payload_addr_block;
  assign Queue_4_1_io_enq_bits_payload_client_xact_id = io_client_acquire_bits_payload_client_xact_id;
  assign Queue_4_1_io_enq_bits_payload_addr_beat = io_client_acquire_bits_payload_addr_beat;
  assign Queue_4_1_io_enq_bits_payload_is_builtin_type = io_client_acquire_bits_payload_is_builtin_type;
  assign Queue_4_1_io_enq_bits_payload_a_type = io_client_acquire_bits_payload_a_type;
  assign Queue_4_1_io_enq_bits_payload_union = io_client_acquire_bits_payload_union;
  assign Queue_4_1_io_enq_bits_payload_data = io_client_acquire_bits_payload_data;
  assign Queue_4_1_io_deq_ready = io_manager_acquire_ready;
  assign Queue_5_1_clk = clk;
  assign Queue_5_1_reset = reset;
  assign Queue_5_1_io_enq_valid = io_manager_probe_valid;
  assign Queue_5_1_io_enq_bits_header_src = io_manager_probe_bits_header_src;
  assign Queue_5_1_io_enq_bits_header_dst = io_manager_probe_bits_header_dst;
  assign Queue_5_1_io_enq_bits_payload_addr_block = io_manager_probe_bits_payload_addr_block;
  assign Queue_5_1_io_enq_bits_payload_p_type = io_manager_probe_bits_payload_p_type;
  assign Queue_5_1_io_deq_ready = io_client_probe_ready;
  assign Queue_6_1_clk = clk;
  assign Queue_6_1_reset = reset;
  assign Queue_6_1_io_enq_valid = io_client_release_valid;
  assign Queue_6_1_io_enq_bits_header_src = io_client_release_bits_header_src;
  assign Queue_6_1_io_enq_bits_header_dst = io_client_release_bits_header_dst;
  assign Queue_6_1_io_enq_bits_payload_addr_beat = io_client_release_bits_payload_addr_beat;
  assign Queue_6_1_io_enq_bits_payload_addr_block = io_client_release_bits_payload_addr_block;
  assign Queue_6_1_io_enq_bits_payload_client_xact_id = io_client_release_bits_payload_client_xact_id;
  assign Queue_6_1_io_enq_bits_payload_voluntary = io_client_release_bits_payload_voluntary;
  assign Queue_6_1_io_enq_bits_payload_r_type = io_client_release_bits_payload_r_type;
  assign Queue_6_1_io_enq_bits_payload_data = io_client_release_bits_payload_data;
  assign Queue_6_1_io_deq_ready = io_manager_release_ready;
  assign Queue_7_1_clk = clk;
  assign Queue_7_1_reset = reset;
  assign Queue_7_1_io_enq_valid = io_manager_grant_valid;
  assign Queue_7_1_io_enq_bits_header_src = io_manager_grant_bits_header_src;
  assign Queue_7_1_io_enq_bits_header_dst = io_manager_grant_bits_header_dst;
  assign Queue_7_1_io_enq_bits_payload_addr_beat = io_manager_grant_bits_payload_addr_beat;
  assign Queue_7_1_io_enq_bits_payload_client_xact_id = io_manager_grant_bits_payload_client_xact_id;
  assign Queue_7_1_io_enq_bits_payload_manager_xact_id = io_manager_grant_bits_payload_manager_xact_id;
  assign Queue_7_1_io_enq_bits_payload_is_builtin_type = io_manager_grant_bits_payload_is_builtin_type;
  assign Queue_7_1_io_enq_bits_payload_g_type = io_manager_grant_bits_payload_g_type;
  assign Queue_7_1_io_enq_bits_payload_data = io_manager_grant_bits_payload_data;
  assign Queue_7_1_io_deq_ready = io_client_grant_ready;
endmodule
module FinishQueue_1(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_manager_xact_id,
  input   io_enq_bits_manager_id,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_manager_xact_id,
  output  io_deq_bits_manager_id,
  output [1:0] io_count
);
  reg [1:0] ram_manager_xact_id [0:1];
  reg [31:0] GEN_0;
  wire [1:0] ram_manager_xact_id_T_264_data;
  wire  ram_manager_xact_id_T_264_addr;
  wire  ram_manager_xact_id_T_264_en;
  wire [1:0] ram_manager_xact_id_T_226_data;
  wire  ram_manager_xact_id_T_226_addr;
  wire  ram_manager_xact_id_T_226_mask;
  wire  ram_manager_xact_id_T_226_en;
  reg  ram_manager_id [0:1];
  reg [31:0] GEN_1;
  wire  ram_manager_id_T_264_data;
  wire  ram_manager_id_T_264_addr;
  wire  ram_manager_id_T_264_en;
  wire  ram_manager_id_T_226_data;
  wire  ram_manager_id_T_226_addr;
  wire  ram_manager_id_T_226_mask;
  wire  ram_manager_id_T_226_en;
  reg  T_218;
  reg [31:0] GEN_2;
  reg  T_220;
  reg [31:0] GEN_3;
  reg  maybe_full;
  reg [31:0] GEN_4;
  wire  ptr_match;
  wire  T_223;
  wire  empty;
  wire  full;
  wire  T_224;
  wire  do_enq;
  wire  T_225;
  wire  do_deq;
  wire [1:0] T_252;
  wire  T_253;
  wire  GEN_7;
  wire [1:0] T_257;
  wire  T_258;
  wire  GEN_8;
  wire  T_259;
  wire  GEN_9;
  wire  T_261;
  wire  T_263;
  wire [1:0] T_287;
  wire  ptr_diff;
  wire  T_288;
  wire [1:0] T_289;
  assign io_enq_ready = T_263;
  assign io_deq_valid = T_261;
  assign io_deq_bits_manager_xact_id = ram_manager_xact_id_T_264_data;
  assign io_deq_bits_manager_id = ram_manager_id_T_264_data;
  assign io_count = T_289;
  assign ram_manager_xact_id_T_264_addr = T_220;
  assign ram_manager_xact_id_T_264_en = 1'h1;
  assign ram_manager_xact_id_T_264_data = ram_manager_xact_id[ram_manager_xact_id_T_264_addr];
  assign ram_manager_xact_id_T_226_data = io_enq_bits_manager_xact_id;
  assign ram_manager_xact_id_T_226_addr = T_218;
  assign ram_manager_xact_id_T_226_mask = do_enq;
  assign ram_manager_xact_id_T_226_en = do_enq;
  assign ram_manager_id_T_264_addr = T_220;
  assign ram_manager_id_T_264_en = 1'h1;
  assign ram_manager_id_T_264_data = ram_manager_id[ram_manager_id_T_264_addr];
  assign ram_manager_id_T_226_data = io_enq_bits_manager_id;
  assign ram_manager_id_T_226_addr = T_218;
  assign ram_manager_id_T_226_mask = do_enq;
  assign ram_manager_id_T_226_en = do_enq;
  assign ptr_match = T_218 == T_220;
  assign T_223 = maybe_full == 1'h0;
  assign empty = ptr_match & T_223;
  assign full = ptr_match & maybe_full;
  assign T_224 = io_enq_ready & io_enq_valid;
  assign do_enq = T_224;
  assign T_225 = io_deq_ready & io_deq_valid;
  assign do_deq = T_225;
  assign T_252 = T_218 + 1'h1;
  assign T_253 = T_252[0:0];
  assign GEN_7 = do_enq ? T_253 : T_218;
  assign T_257 = T_220 + 1'h1;
  assign T_258 = T_257[0:0];
  assign GEN_8 = do_deq ? T_258 : T_220;
  assign T_259 = do_enq != do_deq;
  assign GEN_9 = T_259 ? do_enq : maybe_full;
  assign T_261 = empty == 1'h0;
  assign T_263 = full == 1'h0;
  assign T_287 = T_218 - T_220;
  assign ptr_diff = T_287[0:0];
  assign T_288 = maybe_full & ptr_match;
  assign T_289 = {T_288,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_manager_xact_id[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_manager_id[initvar] = GEN_1[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_2 = {1{$random}};
  T_218 = GEN_2[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_3 = {1{$random}};
  T_220 = GEN_3[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_4 = {1{$random}};
  maybe_full = GEN_4[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_manager_xact_id_T_226_en & ram_manager_xact_id_T_226_mask) begin
      ram_manager_xact_id[ram_manager_xact_id_T_226_addr] <= ram_manager_xact_id_T_226_data;
    end
    if(ram_manager_id_T_226_en & ram_manager_id_T_226_mask) begin
      ram_manager_id[ram_manager_id_T_226_addr] <= ram_manager_id_T_226_data;
    end
    if(reset) begin
      T_218 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_218 <= T_253;
      end
    end
    if(reset) begin
      T_220 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_220 <= T_258;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_259) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module FinishUnit(
  input   clk,
  input   reset,
  output  io_grant_ready,
  input   io_grant_valid,
  input  [1:0] io_grant_bits_header_src,
  input  [1:0] io_grant_bits_header_dst,
  input  [2:0] io_grant_bits_payload_addr_beat,
  input   io_grant_bits_payload_client_xact_id,
  input  [1:0] io_grant_bits_payload_manager_xact_id,
  input   io_grant_bits_payload_is_builtin_type,
  input  [3:0] io_grant_bits_payload_g_type,
  input  [63:0] io_grant_bits_payload_data,
  input   io_refill_ready,
  output  io_refill_valid,
  output [2:0] io_refill_bits_addr_beat,
  output  io_refill_bits_client_xact_id,
  output [1:0] io_refill_bits_manager_xact_id,
  output  io_refill_bits_is_builtin_type,
  output [3:0] io_refill_bits_g_type,
  output [63:0] io_refill_bits_data,
  input   io_finish_ready,
  output  io_finish_valid,
  output [1:0] io_finish_bits_header_src,
  output [1:0] io_finish_bits_header_dst,
  output [1:0] io_finish_bits_payload_manager_xact_id,
  output  io_ready
);
  wire  T_1035;
  wire [2:0] T_1044_0;
  wire [3:0] GEN_1;
  wire  T_1046;
  wire  T_1047;
  wire  T_1048;
  wire  T_1050;
  reg [2:0] T_1052;
  reg [31:0] GEN_3;
  wire  T_1054;
  wire [3:0] T_1056;
  wire [2:0] T_1057;
  wire [2:0] GEN_0;
  wire  T_1058;
  wire  T_1060;
  wire  FinishQueue_1_1_clk;
  wire  FinishQueue_1_1_reset;
  wire  FinishQueue_1_1_io_enq_ready;
  wire  FinishQueue_1_1_io_enq_valid;
  wire [1:0] FinishQueue_1_1_io_enq_bits_manager_xact_id;
  wire  FinishQueue_1_1_io_enq_bits_manager_id;
  wire  FinishQueue_1_1_io_deq_ready;
  wire  FinishQueue_1_1_io_deq_valid;
  wire [1:0] FinishQueue_1_1_io_deq_bits_manager_xact_id;
  wire  FinishQueue_1_1_io_deq_bits_manager_id;
  wire [1:0] FinishQueue_1_1_io_count;
  wire  T_1090;
  wire  T_1092;
  wire  T_1094;
  wire [2:0] T_1102_0;
  wire [3:0] GEN_2;
  wire  T_1104;
  wire  T_1106;
  wire  T_1109;
  wire  T_1110;
  wire  T_1111;
  wire [1:0] T_1134_manager_xact_id;
  wire  T_1167;
  wire  T_1168;
  wire  T_1169;
  wire  T_1182;
  FinishQueue_1 FinishQueue_1_1 (
    .clk(FinishQueue_1_1_clk),
    .reset(FinishQueue_1_1_reset),
    .io_enq_ready(FinishQueue_1_1_io_enq_ready),
    .io_enq_valid(FinishQueue_1_1_io_enq_valid),
    .io_enq_bits_manager_xact_id(FinishQueue_1_1_io_enq_bits_manager_xact_id),
    .io_enq_bits_manager_id(FinishQueue_1_1_io_enq_bits_manager_id),
    .io_deq_ready(FinishQueue_1_1_io_deq_ready),
    .io_deq_valid(FinishQueue_1_1_io_deq_valid),
    .io_deq_bits_manager_xact_id(FinishQueue_1_1_io_deq_bits_manager_xact_id),
    .io_deq_bits_manager_id(FinishQueue_1_1_io_deq_bits_manager_id),
    .io_count(FinishQueue_1_1_io_count)
  );
  assign io_grant_ready = T_1182;
  assign io_refill_valid = T_1169;
  assign io_refill_bits_addr_beat = io_grant_bits_payload_addr_beat;
  assign io_refill_bits_client_xact_id = io_grant_bits_payload_client_xact_id;
  assign io_refill_bits_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign io_refill_bits_is_builtin_type = io_grant_bits_payload_is_builtin_type;
  assign io_refill_bits_g_type = io_grant_bits_payload_g_type;
  assign io_refill_bits_data = io_grant_bits_payload_data;
  assign io_finish_valid = FinishQueue_1_1_io_deq_valid;
  assign io_finish_bits_header_src = 2'h1;
  assign io_finish_bits_header_dst = {{1'd0}, FinishQueue_1_1_io_deq_bits_manager_id};
  assign io_finish_bits_payload_manager_xact_id = FinishQueue_1_1_io_deq_bits_manager_xact_id;
  assign io_ready = FinishQueue_1_1_io_enq_ready;
  assign T_1035 = io_grant_ready & io_grant_valid;
  assign T_1044_0 = 3'h5;
  assign GEN_1 = {{1'd0}, T_1044_0};
  assign T_1046 = io_grant_bits_payload_g_type == GEN_1;
  assign T_1047 = io_grant_bits_payload_g_type == 4'h0;
  assign T_1048 = io_grant_bits_payload_is_builtin_type ? T_1046 : T_1047;
  assign T_1050 = T_1035 & T_1048;
  assign T_1054 = T_1052 == 3'h7;
  assign T_1056 = T_1052 + 3'h1;
  assign T_1057 = T_1056[2:0];
  assign GEN_0 = T_1050 ? T_1057 : T_1052;
  assign T_1058 = T_1050 & T_1054;
  assign T_1060 = T_1048 ? T_1058 : T_1035;
  assign FinishQueue_1_1_clk = clk;
  assign FinishQueue_1_1_reset = reset;
  assign FinishQueue_1_1_io_enq_valid = T_1111;
  assign FinishQueue_1_1_io_enq_bits_manager_xact_id = T_1134_manager_xact_id;
  assign FinishQueue_1_1_io_enq_bits_manager_id = io_grant_bits_header_src[0];
  assign FinishQueue_1_1_io_deq_ready = io_finish_ready;
  assign T_1090 = io_grant_bits_payload_is_builtin_type & T_1047;
  assign T_1092 = T_1090 == 1'h0;
  assign T_1094 = T_1035 & T_1092;
  assign T_1102_0 = 3'h5;
  assign GEN_2 = {{1'd0}, T_1102_0};
  assign T_1104 = io_grant_bits_payload_g_type == GEN_2;
  assign T_1106 = io_grant_bits_payload_is_builtin_type ? T_1104 : T_1047;
  assign T_1109 = T_1106 == 1'h0;
  assign T_1110 = T_1109 | T_1060;
  assign T_1111 = T_1094 & T_1110;
  assign T_1134_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign T_1167 = T_1092 == 1'h0;
  assign T_1168 = FinishQueue_1_1_io_enq_ready | T_1167;
  assign T_1169 = T_1168 & io_grant_valid;
  assign T_1182 = T_1168 & io_refill_ready;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_3 = {1{$random}};
  T_1052 = GEN_3[2:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1052 <= 3'h0;
    end else begin
      if(T_1050) begin
        T_1052 <= T_1057;
      end
    end
  end
endmodule
module ClientUncachedTileLinkNetworkPort(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [25:0] io_client_acquire_bits_addr_block,
  input   io_client_acquire_bits_client_xact_id,
  input  [2:0] io_client_acquire_bits_addr_beat,
  input   io_client_acquire_bits_is_builtin_type,
  input  [2:0] io_client_acquire_bits_a_type,
  input  [11:0] io_client_acquire_bits_union,
  input  [63:0] io_client_acquire_bits_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [2:0] io_client_grant_bits_addr_beat,
  output  io_client_grant_bits_client_xact_id,
  output [1:0] io_client_grant_bits_manager_xact_id,
  output  io_client_grant_bits_is_builtin_type,
  output [3:0] io_client_grant_bits_g_type,
  output [63:0] io_client_grant_bits_data,
  input   io_network_acquire_ready,
  output  io_network_acquire_valid,
  output [1:0] io_network_acquire_bits_header_src,
  output [1:0] io_network_acquire_bits_header_dst,
  output [25:0] io_network_acquire_bits_payload_addr_block,
  output  io_network_acquire_bits_payload_client_xact_id,
  output [2:0] io_network_acquire_bits_payload_addr_beat,
  output  io_network_acquire_bits_payload_is_builtin_type,
  output [2:0] io_network_acquire_bits_payload_a_type,
  output [11:0] io_network_acquire_bits_payload_union,
  output [63:0] io_network_acquire_bits_payload_data,
  output  io_network_grant_ready,
  input   io_network_grant_valid,
  input  [1:0] io_network_grant_bits_header_src,
  input  [1:0] io_network_grant_bits_header_dst,
  input  [2:0] io_network_grant_bits_payload_addr_beat,
  input   io_network_grant_bits_payload_client_xact_id,
  input  [1:0] io_network_grant_bits_payload_manager_xact_id,
  input   io_network_grant_bits_payload_is_builtin_type,
  input  [3:0] io_network_grant_bits_payload_g_type,
  input  [63:0] io_network_grant_bits_payload_data,
  input   io_network_finish_ready,
  output  io_network_finish_valid,
  output [1:0] io_network_finish_bits_header_src,
  output [1:0] io_network_finish_bits_header_dst,
  output [1:0] io_network_finish_bits_payload_manager_xact_id,
  output  io_network_probe_ready,
  input   io_network_probe_valid,
  input  [1:0] io_network_probe_bits_header_src,
  input  [1:0] io_network_probe_bits_header_dst,
  input  [25:0] io_network_probe_bits_payload_addr_block,
  input  [1:0] io_network_probe_bits_payload_p_type,
  input   io_network_release_ready,
  output  io_network_release_valid,
  output [1:0] io_network_release_bits_header_src,
  output [1:0] io_network_release_bits_header_dst,
  output [2:0] io_network_release_bits_payload_addr_beat,
  output [25:0] io_network_release_bits_payload_addr_block,
  output  io_network_release_bits_payload_client_xact_id,
  output  io_network_release_bits_payload_voluntary,
  output [2:0] io_network_release_bits_payload_r_type,
  output [63:0] io_network_release_bits_payload_data
);
  wire  finisher_clk;
  wire  finisher_reset;
  wire  finisher_io_grant_ready;
  wire  finisher_io_grant_valid;
  wire [1:0] finisher_io_grant_bits_header_src;
  wire [1:0] finisher_io_grant_bits_header_dst;
  wire [2:0] finisher_io_grant_bits_payload_addr_beat;
  wire  finisher_io_grant_bits_payload_client_xact_id;
  wire [1:0] finisher_io_grant_bits_payload_manager_xact_id;
  wire  finisher_io_grant_bits_payload_is_builtin_type;
  wire [3:0] finisher_io_grant_bits_payload_g_type;
  wire [63:0] finisher_io_grant_bits_payload_data;
  wire  finisher_io_refill_ready;
  wire  finisher_io_refill_valid;
  wire [2:0] finisher_io_refill_bits_addr_beat;
  wire  finisher_io_refill_bits_client_xact_id;
  wire [1:0] finisher_io_refill_bits_manager_xact_id;
  wire  finisher_io_refill_bits_is_builtin_type;
  wire [3:0] finisher_io_refill_bits_g_type;
  wire [63:0] finisher_io_refill_bits_data;
  wire  finisher_io_finish_ready;
  wire  finisher_io_finish_valid;
  wire [1:0] finisher_io_finish_bits_header_src;
  wire [1:0] finisher_io_finish_bits_header_dst;
  wire [1:0] finisher_io_finish_bits_payload_manager_xact_id;
  wire  finisher_io_ready;
  wire  acq_with_header_ready;
  wire  acq_with_header_valid;
  wire [1:0] acq_with_header_bits_header_src;
  wire [1:0] acq_with_header_bits_header_dst;
  wire [25:0] acq_with_header_bits_payload_addr_block;
  wire  acq_with_header_bits_payload_client_xact_id;
  wire [2:0] acq_with_header_bits_payload_addr_beat;
  wire  acq_with_header_bits_payload_is_builtin_type;
  wire [2:0] acq_with_header_bits_payload_a_type;
  wire [11:0] acq_with_header_bits_payload_union;
  wire [63:0] acq_with_header_bits_payload_data;
  wire [31:0] GEN_0;
  wire [31:0] T_3330;
  wire  T_3332;
  wire  T_3334;
  wire  T_3335;
  wire  T_3338;
  wire  T_3339;
  wire  T_3340;
  reg [1:0] GEN_1;
  reg [31:0] GEN_9;
  reg [1:0] GEN_2;
  reg [31:0] GEN_10;
  reg [2:0] GEN_3;
  reg [31:0] GEN_11;
  reg [25:0] GEN_4;
  reg [31:0] GEN_12;
  reg  GEN_5;
  reg [31:0] GEN_13;
  reg  GEN_6;
  reg [31:0] GEN_14;
  reg [2:0] GEN_7;
  reg [31:0] GEN_15;
  reg [63:0] GEN_8;
  reg [63:0] GEN_16;
  FinishUnit finisher (
    .clk(finisher_clk),
    .reset(finisher_reset),
    .io_grant_ready(finisher_io_grant_ready),
    .io_grant_valid(finisher_io_grant_valid),
    .io_grant_bits_header_src(finisher_io_grant_bits_header_src),
    .io_grant_bits_header_dst(finisher_io_grant_bits_header_dst),
    .io_grant_bits_payload_addr_beat(finisher_io_grant_bits_payload_addr_beat),
    .io_grant_bits_payload_client_xact_id(finisher_io_grant_bits_payload_client_xact_id),
    .io_grant_bits_payload_manager_xact_id(finisher_io_grant_bits_payload_manager_xact_id),
    .io_grant_bits_payload_is_builtin_type(finisher_io_grant_bits_payload_is_builtin_type),
    .io_grant_bits_payload_g_type(finisher_io_grant_bits_payload_g_type),
    .io_grant_bits_payload_data(finisher_io_grant_bits_payload_data),
    .io_refill_ready(finisher_io_refill_ready),
    .io_refill_valid(finisher_io_refill_valid),
    .io_refill_bits_addr_beat(finisher_io_refill_bits_addr_beat),
    .io_refill_bits_client_xact_id(finisher_io_refill_bits_client_xact_id),
    .io_refill_bits_manager_xact_id(finisher_io_refill_bits_manager_xact_id),
    .io_refill_bits_is_builtin_type(finisher_io_refill_bits_is_builtin_type),
    .io_refill_bits_g_type(finisher_io_refill_bits_g_type),
    .io_refill_bits_data(finisher_io_refill_bits_data),
    .io_finish_ready(finisher_io_finish_ready),
    .io_finish_valid(finisher_io_finish_valid),
    .io_finish_bits_header_src(finisher_io_finish_bits_header_src),
    .io_finish_bits_header_dst(finisher_io_finish_bits_header_dst),
    .io_finish_bits_payload_manager_xact_id(finisher_io_finish_bits_payload_manager_xact_id),
    .io_ready(finisher_io_ready)
  );
  assign io_client_acquire_ready = acq_with_header_ready;
  assign io_client_grant_valid = finisher_io_refill_valid;
  assign io_client_grant_bits_addr_beat = finisher_io_refill_bits_addr_beat;
  assign io_client_grant_bits_client_xact_id = finisher_io_refill_bits_client_xact_id;
  assign io_client_grant_bits_manager_xact_id = finisher_io_refill_bits_manager_xact_id;
  assign io_client_grant_bits_is_builtin_type = finisher_io_refill_bits_is_builtin_type;
  assign io_client_grant_bits_g_type = finisher_io_refill_bits_g_type;
  assign io_client_grant_bits_data = finisher_io_refill_bits_data;
  assign io_network_acquire_valid = T_3339;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign io_network_grant_ready = finisher_io_grant_ready;
  assign io_network_finish_valid = finisher_io_finish_valid;
  assign io_network_finish_bits_header_src = finisher_io_finish_bits_header_src;
  assign io_network_finish_bits_header_dst = finisher_io_finish_bits_header_dst;
  assign io_network_finish_bits_payload_manager_xact_id = finisher_io_finish_bits_payload_manager_xact_id;
  assign io_network_probe_ready = 1'h0;
  assign io_network_release_valid = 1'h0;
  assign io_network_release_bits_header_src = GEN_1;
  assign io_network_release_bits_header_dst = GEN_2;
  assign io_network_release_bits_payload_addr_beat = GEN_3;
  assign io_network_release_bits_payload_addr_block = GEN_4;
  assign io_network_release_bits_payload_client_xact_id = GEN_5;
  assign io_network_release_bits_payload_voluntary = GEN_6;
  assign io_network_release_bits_payload_r_type = GEN_7;
  assign io_network_release_bits_payload_data = GEN_8;
  assign finisher_clk = clk;
  assign finisher_reset = reset;
  assign finisher_io_grant_valid = io_network_grant_valid;
  assign finisher_io_grant_bits_header_src = io_network_grant_bits_header_src;
  assign finisher_io_grant_bits_header_dst = io_network_grant_bits_header_dst;
  assign finisher_io_grant_bits_payload_addr_beat = io_network_grant_bits_payload_addr_beat;
  assign finisher_io_grant_bits_payload_client_xact_id = io_network_grant_bits_payload_client_xact_id;
  assign finisher_io_grant_bits_payload_manager_xact_id = io_network_grant_bits_payload_manager_xact_id;
  assign finisher_io_grant_bits_payload_is_builtin_type = io_network_grant_bits_payload_is_builtin_type;
  assign finisher_io_grant_bits_payload_g_type = io_network_grant_bits_payload_g_type;
  assign finisher_io_grant_bits_payload_data = io_network_grant_bits_payload_data;
  assign finisher_io_refill_ready = io_client_grant_ready;
  assign finisher_io_finish_ready = io_network_finish_ready;
  assign acq_with_header_ready = T_3340;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign acq_with_header_bits_header_src = 2'h1;
  assign acq_with_header_bits_header_dst = {{1'd0}, T_3338};
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign GEN_0 = {{6'd0}, io_client_acquire_bits_addr_block};
  assign T_3330 = GEN_0 << 6;
  assign T_3332 = 32'h80000000 <= T_3330;
  assign T_3334 = T_3330 < 32'h90000000;
  assign T_3335 = T_3332 & T_3334;
  assign T_3338 = T_3335 ? 1'h0 : 1'h1;
  assign T_3339 = acq_with_header_valid & finisher_io_ready;
  assign T_3340 = io_network_acquire_ready & finisher_io_ready;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_9 = {1{$random}};
  GEN_1 = GEN_9[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_10 = {1{$random}};
  GEN_2 = GEN_10[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_11 = {1{$random}};
  GEN_3 = GEN_11[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_12 = {1{$random}};
  GEN_4 = GEN_12[25:0];
  `endif
  `ifdef RANDOMIZE
  GEN_13 = {1{$random}};
  GEN_5 = GEN_13[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_14 = {1{$random}};
  GEN_6 = GEN_14[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_15 = {1{$random}};
  GEN_7 = GEN_15[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_16 = {2{$random}};
  GEN_8 = GEN_16[63:0];
  `endif
  end
`endif
endmodule
module ManagerTileLinkNetworkPort(
  input   clk,
  input   reset,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [25:0] io_manager_acquire_bits_addr_block,
  output  io_manager_acquire_bits_client_xact_id,
  output [2:0] io_manager_acquire_bits_addr_beat,
  output  io_manager_acquire_bits_is_builtin_type,
  output [2:0] io_manager_acquire_bits_a_type,
  output [11:0] io_manager_acquire_bits_union,
  output [63:0] io_manager_acquire_bits_data,
  output  io_manager_acquire_bits_client_id,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [2:0] io_manager_grant_bits_addr_beat,
  input   io_manager_grant_bits_client_xact_id,
  input  [1:0] io_manager_grant_bits_manager_xact_id,
  input   io_manager_grant_bits_is_builtin_type,
  input  [3:0] io_manager_grant_bits_g_type,
  input  [63:0] io_manager_grant_bits_data,
  input   io_manager_grant_bits_client_id,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [1:0] io_manager_finish_bits_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [25:0] io_manager_probe_bits_addr_block,
  input  [1:0] io_manager_probe_bits_p_type,
  input   io_manager_probe_bits_client_id,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [2:0] io_manager_release_bits_addr_beat,
  output [25:0] io_manager_release_bits_addr_block,
  output  io_manager_release_bits_client_xact_id,
  output  io_manager_release_bits_voluntary,
  output [2:0] io_manager_release_bits_r_type,
  output [63:0] io_manager_release_bits_data,
  output  io_manager_release_bits_client_id,
  output  io_network_acquire_ready,
  input   io_network_acquire_valid,
  input  [1:0] io_network_acquire_bits_header_src,
  input  [1:0] io_network_acquire_bits_header_dst,
  input  [25:0] io_network_acquire_bits_payload_addr_block,
  input   io_network_acquire_bits_payload_client_xact_id,
  input  [2:0] io_network_acquire_bits_payload_addr_beat,
  input   io_network_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_network_acquire_bits_payload_a_type,
  input  [11:0] io_network_acquire_bits_payload_union,
  input  [63:0] io_network_acquire_bits_payload_data,
  input   io_network_grant_ready,
  output  io_network_grant_valid,
  output [1:0] io_network_grant_bits_header_src,
  output [1:0] io_network_grant_bits_header_dst,
  output [2:0] io_network_grant_bits_payload_addr_beat,
  output  io_network_grant_bits_payload_client_xact_id,
  output [1:0] io_network_grant_bits_payload_manager_xact_id,
  output  io_network_grant_bits_payload_is_builtin_type,
  output [3:0] io_network_grant_bits_payload_g_type,
  output [63:0] io_network_grant_bits_payload_data,
  output  io_network_finish_ready,
  input   io_network_finish_valid,
  input  [1:0] io_network_finish_bits_header_src,
  input  [1:0] io_network_finish_bits_header_dst,
  input  [1:0] io_network_finish_bits_payload_manager_xact_id,
  input   io_network_probe_ready,
  output  io_network_probe_valid,
  output [1:0] io_network_probe_bits_header_src,
  output [1:0] io_network_probe_bits_header_dst,
  output [25:0] io_network_probe_bits_payload_addr_block,
  output [1:0] io_network_probe_bits_payload_p_type,
  output  io_network_release_ready,
  input   io_network_release_valid,
  input  [1:0] io_network_release_bits_header_src,
  input  [1:0] io_network_release_bits_header_dst,
  input  [2:0] io_network_release_bits_payload_addr_beat,
  input  [25:0] io_network_release_bits_payload_addr_block,
  input   io_network_release_bits_payload_client_xact_id,
  input   io_network_release_bits_payload_voluntary,
  input  [2:0] io_network_release_bits_payload_r_type,
  input  [63:0] io_network_release_bits_payload_data
);
  wire  T_6043_ready;
  wire  T_6043_valid;
  wire [1:0] T_6043_bits_header_src;
  wire [1:0] T_6043_bits_header_dst;
  wire [2:0] T_6043_bits_payload_addr_beat;
  wire  T_6043_bits_payload_client_xact_id;
  wire [1:0] T_6043_bits_payload_manager_xact_id;
  wire  T_6043_bits_payload_is_builtin_type;
  wire [3:0] T_6043_bits_payload_g_type;
  wire [63:0] T_6043_bits_payload_data;
  wire  T_6043_bits_payload_client_id;
  wire  T_6598_ready;
  wire  T_6598_valid;
  wire [1:0] T_6598_bits_header_src;
  wire [1:0] T_6598_bits_header_dst;
  wire [25:0] T_6598_bits_payload_addr_block;
  wire [1:0] T_6598_bits_payload_p_type;
  wire  T_6598_bits_payload_client_id;
  wire  T_6877_ready;
  wire  T_6877_valid;
  wire [25:0] T_6877_bits_addr_block;
  wire  T_6877_bits_client_xact_id;
  wire [2:0] T_6877_bits_addr_beat;
  wire  T_6877_bits_is_builtin_type;
  wire [2:0] T_6877_bits_a_type;
  wire [11:0] T_6877_bits_union;
  wire [63:0] T_6877_bits_data;
  wire  T_6993_ready;
  wire  T_6993_valid;
  wire [2:0] T_6993_bits_addr_beat;
  wire [25:0] T_6993_bits_addr_block;
  wire  T_6993_bits_client_xact_id;
  wire  T_6993_bits_voluntary;
  wire [2:0] T_6993_bits_r_type;
  wire [63:0] T_6993_bits_data;
  wire  T_7097_ready;
  wire  T_7097_valid;
  wire [1:0] T_7097_bits_manager_xact_id;
  assign io_manager_acquire_valid = T_6877_valid;
  assign io_manager_acquire_bits_addr_block = T_6877_bits_addr_block;
  assign io_manager_acquire_bits_client_xact_id = T_6877_bits_client_xact_id;
  assign io_manager_acquire_bits_addr_beat = T_6877_bits_addr_beat;
  assign io_manager_acquire_bits_is_builtin_type = T_6877_bits_is_builtin_type;
  assign io_manager_acquire_bits_a_type = T_6877_bits_a_type;
  assign io_manager_acquire_bits_union = T_6877_bits_union;
  assign io_manager_acquire_bits_data = T_6877_bits_data;
  assign io_manager_acquire_bits_client_id = io_network_acquire_bits_header_src[0];
  assign io_manager_grant_ready = T_6043_ready;
  assign io_manager_finish_valid = T_7097_valid;
  assign io_manager_finish_bits_manager_xact_id = T_7097_bits_manager_xact_id;
  assign io_manager_probe_ready = T_6598_ready;
  assign io_manager_release_valid = T_6993_valid;
  assign io_manager_release_bits_addr_beat = T_6993_bits_addr_beat;
  assign io_manager_release_bits_addr_block = T_6993_bits_addr_block;
  assign io_manager_release_bits_client_xact_id = T_6993_bits_client_xact_id;
  assign io_manager_release_bits_voluntary = T_6993_bits_voluntary;
  assign io_manager_release_bits_r_type = T_6993_bits_r_type;
  assign io_manager_release_bits_data = T_6993_bits_data;
  assign io_manager_release_bits_client_id = io_network_release_bits_header_src[0];
  assign io_network_acquire_ready = T_6877_ready;
  assign io_network_grant_valid = T_6043_valid;
  assign io_network_grant_bits_header_src = T_6043_bits_header_src;
  assign io_network_grant_bits_header_dst = T_6043_bits_header_dst;
  assign io_network_grant_bits_payload_addr_beat = T_6043_bits_payload_addr_beat;
  assign io_network_grant_bits_payload_client_xact_id = T_6043_bits_payload_client_xact_id;
  assign io_network_grant_bits_payload_manager_xact_id = T_6043_bits_payload_manager_xact_id;
  assign io_network_grant_bits_payload_is_builtin_type = T_6043_bits_payload_is_builtin_type;
  assign io_network_grant_bits_payload_g_type = T_6043_bits_payload_g_type;
  assign io_network_grant_bits_payload_data = T_6043_bits_payload_data;
  assign io_network_finish_ready = T_7097_ready;
  assign io_network_probe_valid = T_6598_valid;
  assign io_network_probe_bits_header_src = T_6598_bits_header_src;
  assign io_network_probe_bits_header_dst = T_6598_bits_header_dst;
  assign io_network_probe_bits_payload_addr_block = T_6598_bits_payload_addr_block;
  assign io_network_probe_bits_payload_p_type = T_6598_bits_payload_p_type;
  assign io_network_release_ready = T_6993_ready;
  assign T_6043_ready = io_network_grant_ready;
  assign T_6043_valid = io_manager_grant_valid;
  assign T_6043_bits_header_src = 2'h0;
  assign T_6043_bits_header_dst = {{1'd0}, io_manager_grant_bits_client_id};
  assign T_6043_bits_payload_addr_beat = io_manager_grant_bits_addr_beat;
  assign T_6043_bits_payload_client_xact_id = io_manager_grant_bits_client_xact_id;
  assign T_6043_bits_payload_manager_xact_id = io_manager_grant_bits_manager_xact_id;
  assign T_6043_bits_payload_is_builtin_type = io_manager_grant_bits_is_builtin_type;
  assign T_6043_bits_payload_g_type = io_manager_grant_bits_g_type;
  assign T_6043_bits_payload_data = io_manager_grant_bits_data;
  assign T_6043_bits_payload_client_id = io_manager_grant_bits_client_id;
  assign T_6598_ready = io_network_probe_ready;
  assign T_6598_valid = io_manager_probe_valid;
  assign T_6598_bits_header_src = 2'h0;
  assign T_6598_bits_header_dst = {{1'd0}, io_manager_probe_bits_client_id};
  assign T_6598_bits_payload_addr_block = io_manager_probe_bits_addr_block;
  assign T_6598_bits_payload_p_type = io_manager_probe_bits_p_type;
  assign T_6598_bits_payload_client_id = io_manager_probe_bits_client_id;
  assign T_6877_ready = io_manager_acquire_ready;
  assign T_6877_valid = io_network_acquire_valid;
  assign T_6877_bits_addr_block = io_network_acquire_bits_payload_addr_block;
  assign T_6877_bits_client_xact_id = io_network_acquire_bits_payload_client_xact_id;
  assign T_6877_bits_addr_beat = io_network_acquire_bits_payload_addr_beat;
  assign T_6877_bits_is_builtin_type = io_network_acquire_bits_payload_is_builtin_type;
  assign T_6877_bits_a_type = io_network_acquire_bits_payload_a_type;
  assign T_6877_bits_union = io_network_acquire_bits_payload_union;
  assign T_6877_bits_data = io_network_acquire_bits_payload_data;
  assign T_6993_ready = io_manager_release_ready;
  assign T_6993_valid = io_network_release_valid;
  assign T_6993_bits_addr_beat = io_network_release_bits_payload_addr_beat;
  assign T_6993_bits_addr_block = io_network_release_bits_payload_addr_block;
  assign T_6993_bits_client_xact_id = io_network_release_bits_payload_client_xact_id;
  assign T_6993_bits_voluntary = io_network_release_bits_payload_voluntary;
  assign T_6993_bits_r_type = io_network_release_bits_payload_r_type;
  assign T_6993_bits_data = io_network_release_bits_payload_data;
  assign T_7097_ready = io_manager_finish_ready;
  assign T_7097_valid = io_network_finish_valid;
  assign T_7097_bits_manager_xact_id = io_network_finish_bits_payload_manager_xact_id;
endmodule
module TileLinkEnqueuer_2(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [1:0] io_client_acquire_bits_header_src,
  input  [1:0] io_client_acquire_bits_header_dst,
  input  [25:0] io_client_acquire_bits_payload_addr_block,
  input   io_client_acquire_bits_payload_client_xact_id,
  input  [2:0] io_client_acquire_bits_payload_addr_beat,
  input   io_client_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_client_acquire_bits_payload_a_type,
  input  [11:0] io_client_acquire_bits_payload_union,
  input  [63:0] io_client_acquire_bits_payload_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [1:0] io_client_grant_bits_header_src,
  output [1:0] io_client_grant_bits_header_dst,
  output [2:0] io_client_grant_bits_payload_addr_beat,
  output  io_client_grant_bits_payload_client_xact_id,
  output [1:0] io_client_grant_bits_payload_manager_xact_id,
  output  io_client_grant_bits_payload_is_builtin_type,
  output [3:0] io_client_grant_bits_payload_g_type,
  output [63:0] io_client_grant_bits_payload_data,
  output  io_client_finish_ready,
  input   io_client_finish_valid,
  input  [1:0] io_client_finish_bits_header_src,
  input  [1:0] io_client_finish_bits_header_dst,
  input  [1:0] io_client_finish_bits_payload_manager_xact_id,
  input   io_client_probe_ready,
  output  io_client_probe_valid,
  output [1:0] io_client_probe_bits_header_src,
  output [1:0] io_client_probe_bits_header_dst,
  output [25:0] io_client_probe_bits_payload_addr_block,
  output [1:0] io_client_probe_bits_payload_p_type,
  output  io_client_release_ready,
  input   io_client_release_valid,
  input  [1:0] io_client_release_bits_header_src,
  input  [1:0] io_client_release_bits_header_dst,
  input  [2:0] io_client_release_bits_payload_addr_beat,
  input  [25:0] io_client_release_bits_payload_addr_block,
  input   io_client_release_bits_payload_client_xact_id,
  input   io_client_release_bits_payload_voluntary,
  input  [2:0] io_client_release_bits_payload_r_type,
  input  [63:0] io_client_release_bits_payload_data,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [1:0] io_manager_acquire_bits_header_src,
  output [1:0] io_manager_acquire_bits_header_dst,
  output [25:0] io_manager_acquire_bits_payload_addr_block,
  output  io_manager_acquire_bits_payload_client_xact_id,
  output [2:0] io_manager_acquire_bits_payload_addr_beat,
  output  io_manager_acquire_bits_payload_is_builtin_type,
  output [2:0] io_manager_acquire_bits_payload_a_type,
  output [11:0] io_manager_acquire_bits_payload_union,
  output [63:0] io_manager_acquire_bits_payload_data,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [1:0] io_manager_grant_bits_header_src,
  input  [1:0] io_manager_grant_bits_header_dst,
  input  [2:0] io_manager_grant_bits_payload_addr_beat,
  input   io_manager_grant_bits_payload_client_xact_id,
  input  [1:0] io_manager_grant_bits_payload_manager_xact_id,
  input   io_manager_grant_bits_payload_is_builtin_type,
  input  [3:0] io_manager_grant_bits_payload_g_type,
  input  [63:0] io_manager_grant_bits_payload_data,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [1:0] io_manager_finish_bits_header_src,
  output [1:0] io_manager_finish_bits_header_dst,
  output [1:0] io_manager_finish_bits_payload_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [1:0] io_manager_probe_bits_header_src,
  input  [1:0] io_manager_probe_bits_header_dst,
  input  [25:0] io_manager_probe_bits_payload_addr_block,
  input  [1:0] io_manager_probe_bits_payload_p_type,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [1:0] io_manager_release_bits_header_src,
  output [1:0] io_manager_release_bits_header_dst,
  output [2:0] io_manager_release_bits_payload_addr_beat,
  output [25:0] io_manager_release_bits_payload_addr_block,
  output  io_manager_release_bits_payload_client_xact_id,
  output  io_manager_release_bits_payload_voluntary,
  output [2:0] io_manager_release_bits_payload_r_type,
  output [63:0] io_manager_release_bits_payload_data
);
  assign io_client_acquire_ready = io_manager_acquire_ready;
  assign io_client_grant_valid = io_manager_grant_valid;
  assign io_client_grant_bits_header_src = io_manager_grant_bits_header_src;
  assign io_client_grant_bits_header_dst = io_manager_grant_bits_header_dst;
  assign io_client_grant_bits_payload_addr_beat = io_manager_grant_bits_payload_addr_beat;
  assign io_client_grant_bits_payload_client_xact_id = io_manager_grant_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_manager_xact_id = io_manager_grant_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_is_builtin_type = io_manager_grant_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_g_type = io_manager_grant_bits_payload_g_type;
  assign io_client_grant_bits_payload_data = io_manager_grant_bits_payload_data;
  assign io_client_finish_ready = io_manager_finish_ready;
  assign io_client_probe_valid = io_manager_probe_valid;
  assign io_client_probe_bits_header_src = io_manager_probe_bits_header_src;
  assign io_client_probe_bits_header_dst = io_manager_probe_bits_header_dst;
  assign io_client_probe_bits_payload_addr_block = io_manager_probe_bits_payload_addr_block;
  assign io_client_probe_bits_payload_p_type = io_manager_probe_bits_payload_p_type;
  assign io_client_release_ready = io_manager_release_ready;
  assign io_manager_acquire_valid = io_client_acquire_valid;
  assign io_manager_acquire_bits_header_src = io_client_acquire_bits_header_src;
  assign io_manager_acquire_bits_header_dst = io_client_acquire_bits_header_dst;
  assign io_manager_acquire_bits_payload_addr_block = io_client_acquire_bits_payload_addr_block;
  assign io_manager_acquire_bits_payload_client_xact_id = io_client_acquire_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_beat = io_client_acquire_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_is_builtin_type = io_client_acquire_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_a_type = io_client_acquire_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_union = io_client_acquire_bits_payload_union;
  assign io_manager_acquire_bits_payload_data = io_client_acquire_bits_payload_data;
  assign io_manager_grant_ready = io_client_grant_ready;
  assign io_manager_finish_valid = io_client_finish_valid;
  assign io_manager_finish_bits_header_src = io_client_finish_bits_header_src;
  assign io_manager_finish_bits_header_dst = io_client_finish_bits_header_dst;
  assign io_manager_finish_bits_payload_manager_xact_id = io_client_finish_bits_payload_manager_xact_id;
  assign io_manager_probe_ready = io_client_probe_ready;
  assign io_manager_release_valid = io_client_release_valid;
  assign io_manager_release_bits_header_src = io_client_release_bits_header_src;
  assign io_manager_release_bits_header_dst = io_client_release_bits_header_dst;
  assign io_manager_release_bits_payload_addr_beat = io_client_release_bits_payload_addr_beat;
  assign io_manager_release_bits_payload_addr_block = io_client_release_bits_payload_addr_block;
  assign io_manager_release_bits_payload_client_xact_id = io_client_release_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_voluntary = io_client_release_bits_payload_voluntary;
  assign io_manager_release_bits_payload_r_type = io_client_release_bits_payload_r_type;
  assign io_manager_release_bits_payload_data = io_client_release_bits_payload_data;
endmodule
module ManagerTileLinkNetworkPort_1(
  input   clk,
  input   reset,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [25:0] io_manager_acquire_bits_addr_block,
  output  io_manager_acquire_bits_client_xact_id,
  output [2:0] io_manager_acquire_bits_addr_beat,
  output  io_manager_acquire_bits_is_builtin_type,
  output [2:0] io_manager_acquire_bits_a_type,
  output [11:0] io_manager_acquire_bits_union,
  output [63:0] io_manager_acquire_bits_data,
  output  io_manager_acquire_bits_client_id,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [2:0] io_manager_grant_bits_addr_beat,
  input   io_manager_grant_bits_client_xact_id,
  input  [1:0] io_manager_grant_bits_manager_xact_id,
  input   io_manager_grant_bits_is_builtin_type,
  input  [3:0] io_manager_grant_bits_g_type,
  input  [63:0] io_manager_grant_bits_data,
  input   io_manager_grant_bits_client_id,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [1:0] io_manager_finish_bits_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [25:0] io_manager_probe_bits_addr_block,
  input  [1:0] io_manager_probe_bits_p_type,
  input   io_manager_probe_bits_client_id,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [2:0] io_manager_release_bits_addr_beat,
  output [25:0] io_manager_release_bits_addr_block,
  output  io_manager_release_bits_client_xact_id,
  output  io_manager_release_bits_voluntary,
  output [2:0] io_manager_release_bits_r_type,
  output [63:0] io_manager_release_bits_data,
  output  io_manager_release_bits_client_id,
  output  io_network_acquire_ready,
  input   io_network_acquire_valid,
  input  [1:0] io_network_acquire_bits_header_src,
  input  [1:0] io_network_acquire_bits_header_dst,
  input  [25:0] io_network_acquire_bits_payload_addr_block,
  input   io_network_acquire_bits_payload_client_xact_id,
  input  [2:0] io_network_acquire_bits_payload_addr_beat,
  input   io_network_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_network_acquire_bits_payload_a_type,
  input  [11:0] io_network_acquire_bits_payload_union,
  input  [63:0] io_network_acquire_bits_payload_data,
  input   io_network_grant_ready,
  output  io_network_grant_valid,
  output [1:0] io_network_grant_bits_header_src,
  output [1:0] io_network_grant_bits_header_dst,
  output [2:0] io_network_grant_bits_payload_addr_beat,
  output  io_network_grant_bits_payload_client_xact_id,
  output [1:0] io_network_grant_bits_payload_manager_xact_id,
  output  io_network_grant_bits_payload_is_builtin_type,
  output [3:0] io_network_grant_bits_payload_g_type,
  output [63:0] io_network_grant_bits_payload_data,
  output  io_network_finish_ready,
  input   io_network_finish_valid,
  input  [1:0] io_network_finish_bits_header_src,
  input  [1:0] io_network_finish_bits_header_dst,
  input  [1:0] io_network_finish_bits_payload_manager_xact_id,
  input   io_network_probe_ready,
  output  io_network_probe_valid,
  output [1:0] io_network_probe_bits_header_src,
  output [1:0] io_network_probe_bits_header_dst,
  output [25:0] io_network_probe_bits_payload_addr_block,
  output [1:0] io_network_probe_bits_payload_p_type,
  output  io_network_release_ready,
  input   io_network_release_valid,
  input  [1:0] io_network_release_bits_header_src,
  input  [1:0] io_network_release_bits_header_dst,
  input  [2:0] io_network_release_bits_payload_addr_beat,
  input  [25:0] io_network_release_bits_payload_addr_block,
  input   io_network_release_bits_payload_client_xact_id,
  input   io_network_release_bits_payload_voluntary,
  input  [2:0] io_network_release_bits_payload_r_type,
  input  [63:0] io_network_release_bits_payload_data
);
  wire  T_6043_ready;
  wire  T_6043_valid;
  wire [1:0] T_6043_bits_header_src;
  wire [1:0] T_6043_bits_header_dst;
  wire [2:0] T_6043_bits_payload_addr_beat;
  wire  T_6043_bits_payload_client_xact_id;
  wire [1:0] T_6043_bits_payload_manager_xact_id;
  wire  T_6043_bits_payload_is_builtin_type;
  wire [3:0] T_6043_bits_payload_g_type;
  wire [63:0] T_6043_bits_payload_data;
  wire  T_6043_bits_payload_client_id;
  wire  T_6598_ready;
  wire  T_6598_valid;
  wire [1:0] T_6598_bits_header_src;
  wire [1:0] T_6598_bits_header_dst;
  wire [25:0] T_6598_bits_payload_addr_block;
  wire [1:0] T_6598_bits_payload_p_type;
  wire  T_6598_bits_payload_client_id;
  wire  T_6877_ready;
  wire  T_6877_valid;
  wire [25:0] T_6877_bits_addr_block;
  wire  T_6877_bits_client_xact_id;
  wire [2:0] T_6877_bits_addr_beat;
  wire  T_6877_bits_is_builtin_type;
  wire [2:0] T_6877_bits_a_type;
  wire [11:0] T_6877_bits_union;
  wire [63:0] T_6877_bits_data;
  wire  T_6993_ready;
  wire  T_6993_valid;
  wire [2:0] T_6993_bits_addr_beat;
  wire [25:0] T_6993_bits_addr_block;
  wire  T_6993_bits_client_xact_id;
  wire  T_6993_bits_voluntary;
  wire [2:0] T_6993_bits_r_type;
  wire [63:0] T_6993_bits_data;
  wire  T_7097_ready;
  wire  T_7097_valid;
  wire [1:0] T_7097_bits_manager_xact_id;
  assign io_manager_acquire_valid = T_6877_valid;
  assign io_manager_acquire_bits_addr_block = T_6877_bits_addr_block;
  assign io_manager_acquire_bits_client_xact_id = T_6877_bits_client_xact_id;
  assign io_manager_acquire_bits_addr_beat = T_6877_bits_addr_beat;
  assign io_manager_acquire_bits_is_builtin_type = T_6877_bits_is_builtin_type;
  assign io_manager_acquire_bits_a_type = T_6877_bits_a_type;
  assign io_manager_acquire_bits_union = T_6877_bits_union;
  assign io_manager_acquire_bits_data = T_6877_bits_data;
  assign io_manager_acquire_bits_client_id = io_network_acquire_bits_header_src[0];
  assign io_manager_grant_ready = T_6043_ready;
  assign io_manager_finish_valid = T_7097_valid;
  assign io_manager_finish_bits_manager_xact_id = T_7097_bits_manager_xact_id;
  assign io_manager_probe_ready = T_6598_ready;
  assign io_manager_release_valid = T_6993_valid;
  assign io_manager_release_bits_addr_beat = T_6993_bits_addr_beat;
  assign io_manager_release_bits_addr_block = T_6993_bits_addr_block;
  assign io_manager_release_bits_client_xact_id = T_6993_bits_client_xact_id;
  assign io_manager_release_bits_voluntary = T_6993_bits_voluntary;
  assign io_manager_release_bits_r_type = T_6993_bits_r_type;
  assign io_manager_release_bits_data = T_6993_bits_data;
  assign io_manager_release_bits_client_id = io_network_release_bits_header_src[0];
  assign io_network_acquire_ready = T_6877_ready;
  assign io_network_grant_valid = T_6043_valid;
  assign io_network_grant_bits_header_src = T_6043_bits_header_src;
  assign io_network_grant_bits_header_dst = T_6043_bits_header_dst;
  assign io_network_grant_bits_payload_addr_beat = T_6043_bits_payload_addr_beat;
  assign io_network_grant_bits_payload_client_xact_id = T_6043_bits_payload_client_xact_id;
  assign io_network_grant_bits_payload_manager_xact_id = T_6043_bits_payload_manager_xact_id;
  assign io_network_grant_bits_payload_is_builtin_type = T_6043_bits_payload_is_builtin_type;
  assign io_network_grant_bits_payload_g_type = T_6043_bits_payload_g_type;
  assign io_network_grant_bits_payload_data = T_6043_bits_payload_data;
  assign io_network_finish_ready = T_7097_ready;
  assign io_network_probe_valid = T_6598_valid;
  assign io_network_probe_bits_header_src = T_6598_bits_header_src;
  assign io_network_probe_bits_header_dst = T_6598_bits_header_dst;
  assign io_network_probe_bits_payload_addr_block = T_6598_bits_payload_addr_block;
  assign io_network_probe_bits_payload_p_type = T_6598_bits_payload_p_type;
  assign io_network_release_ready = T_6993_ready;
  assign T_6043_ready = io_network_grant_ready;
  assign T_6043_valid = io_manager_grant_valid;
  assign T_6043_bits_header_src = 2'h1;
  assign T_6043_bits_header_dst = {{1'd0}, io_manager_grant_bits_client_id};
  assign T_6043_bits_payload_addr_beat = io_manager_grant_bits_addr_beat;
  assign T_6043_bits_payload_client_xact_id = io_manager_grant_bits_client_xact_id;
  assign T_6043_bits_payload_manager_xact_id = io_manager_grant_bits_manager_xact_id;
  assign T_6043_bits_payload_is_builtin_type = io_manager_grant_bits_is_builtin_type;
  assign T_6043_bits_payload_g_type = io_manager_grant_bits_g_type;
  assign T_6043_bits_payload_data = io_manager_grant_bits_data;
  assign T_6043_bits_payload_client_id = io_manager_grant_bits_client_id;
  assign T_6598_ready = io_network_probe_ready;
  assign T_6598_valid = io_manager_probe_valid;
  assign T_6598_bits_header_src = 2'h1;
  assign T_6598_bits_header_dst = {{1'd0}, io_manager_probe_bits_client_id};
  assign T_6598_bits_payload_addr_block = io_manager_probe_bits_addr_block;
  assign T_6598_bits_payload_p_type = io_manager_probe_bits_p_type;
  assign T_6598_bits_payload_client_id = io_manager_probe_bits_client_id;
  assign T_6877_ready = io_manager_acquire_ready;
  assign T_6877_valid = io_network_acquire_valid;
  assign T_6877_bits_addr_block = io_network_acquire_bits_payload_addr_block;
  assign T_6877_bits_client_xact_id = io_network_acquire_bits_payload_client_xact_id;
  assign T_6877_bits_addr_beat = io_network_acquire_bits_payload_addr_beat;
  assign T_6877_bits_is_builtin_type = io_network_acquire_bits_payload_is_builtin_type;
  assign T_6877_bits_a_type = io_network_acquire_bits_payload_a_type;
  assign T_6877_bits_union = io_network_acquire_bits_payload_union;
  assign T_6877_bits_data = io_network_acquire_bits_payload_data;
  assign T_6993_ready = io_manager_release_ready;
  assign T_6993_valid = io_network_release_valid;
  assign T_6993_bits_addr_beat = io_network_release_bits_payload_addr_beat;
  assign T_6993_bits_addr_block = io_network_release_bits_payload_addr_block;
  assign T_6993_bits_client_xact_id = io_network_release_bits_payload_client_xact_id;
  assign T_6993_bits_voluntary = io_network_release_bits_payload_voluntary;
  assign T_6993_bits_r_type = io_network_release_bits_payload_r_type;
  assign T_6993_bits_data = io_network_release_bits_payload_data;
  assign T_7097_ready = io_manager_finish_ready;
  assign T_7097_valid = io_network_finish_valid;
  assign T_7097_bits_manager_xact_id = io_network_finish_bits_payload_manager_xact_id;
endmodule
module LockingRRArbiter(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input   io_in_0_bits_payload_client_xact_id,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input   io_in_0_bits_payload_is_builtin_type,
  input  [2:0] io_in_0_bits_payload_a_type,
  input  [11:0] io_in_0_bits_payload_union,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input   io_in_1_bits_payload_client_xact_id,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input   io_in_1_bits_payload_is_builtin_type,
  input  [2:0] io_in_1_bits_payload_a_type,
  input  [11:0] io_in_1_bits_payload_union,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input   io_in_2_bits_payload_client_xact_id,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input   io_in_2_bits_payload_is_builtin_type,
  input  [2:0] io_in_2_bits_payload_a_type,
  input  [11:0] io_in_2_bits_payload_union,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input   io_in_3_bits_payload_client_xact_id,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input   io_in_3_bits_payload_is_builtin_type,
  input  [2:0] io_in_3_bits_payload_a_type,
  input  [11:0] io_in_3_bits_payload_union,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_ready,
  output  io_out_valid,
  output [1:0] io_out_bits_header_src,
  output [1:0] io_out_bits_header_dst,
  output [25:0] io_out_bits_payload_addr_block,
  output  io_out_bits_payload_client_xact_id,
  output [2:0] io_out_bits_payload_addr_beat,
  output  io_out_bits_payload_is_builtin_type,
  output [2:0] io_out_bits_payload_a_type,
  output [11:0] io_out_bits_payload_union,
  output [63:0] io_out_bits_payload_data,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire [1:0] GEN_1;
  wire [1:0] GEN_13;
  wire [1:0] GEN_14;
  wire [1:0] GEN_15;
  wire [1:0] GEN_2;
  wire [1:0] GEN_16;
  wire [1:0] GEN_17;
  wire [1:0] GEN_18;
  wire [25:0] GEN_3;
  wire [25:0] GEN_19;
  wire [25:0] GEN_20;
  wire [25:0] GEN_21;
  wire  GEN_4;
  wire  GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire [2:0] GEN_5;
  wire [2:0] GEN_25;
  wire [2:0] GEN_26;
  wire [2:0] GEN_27;
  wire  GEN_6;
  wire  GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire [2:0] GEN_7;
  wire [2:0] GEN_31;
  wire [2:0] GEN_32;
  wire [2:0] GEN_33;
  wire [11:0] GEN_8;
  wire [11:0] GEN_34;
  wire [11:0] GEN_35;
  wire [11:0] GEN_36;
  wire [63:0] GEN_9;
  wire [63:0] GEN_37;
  wire [63:0] GEN_38;
  wire [63:0] GEN_39;
  reg [2:0] T_1134;
  reg [31:0] GEN_50;
  reg [1:0] T_1136;
  reg [31:0] GEN_51;
  wire  T_1138;
  wire [2:0] T_1147_0;
  wire  T_1149;
  wire  T_1150;
  wire  T_1151;
  wire  T_1152;
  wire [3:0] T_1156;
  wire [2:0] T_1157;
  wire [1:0] GEN_40;
  wire [2:0] GEN_41;
  wire [1:0] GEN_42;
  reg [1:0] lastGrant;
  reg [31:0] GEN_52;
  wire [1:0] GEN_43;
  wire  T_1162;
  wire  T_1164;
  wire  T_1166;
  wire  T_1168;
  wire  T_1169;
  wire  T_1170;
  wire  T_1173;
  wire  T_1174;
  wire  T_1175;
  wire  T_1176;
  wire  T_1177;
  wire  T_1181;
  wire  T_1183;
  wire  T_1185;
  wire  T_1187;
  wire  T_1189;
  wire  T_1191;
  wire  T_1195;
  wire  T_1196;
  wire  T_1197;
  wire  T_1198;
  wire  T_1199;
  wire  T_1201;
  wire  T_1202;
  wire  T_1203;
  wire  T_1205;
  wire  T_1206;
  wire  T_1207;
  wire  T_1209;
  wire  T_1210;
  wire  T_1211;
  wire  T_1213;
  wire  T_1214;
  wire  T_1215;
  wire [1:0] GEN_44;
  wire [1:0] GEN_45;
  wire [1:0] GEN_46;
  wire [1:0] GEN_47;
  wire [1:0] GEN_48;
  wire [1:0] GEN_49;
  assign io_in_0_ready = T_1203;
  assign io_in_1_ready = T_1207;
  assign io_in_2_ready = T_1211;
  assign io_in_3_ready = T_1215;
  assign io_out_valid = GEN_0;
  assign io_out_bits_header_src = GEN_1;
  assign io_out_bits_header_dst = GEN_2;
  assign io_out_bits_payload_addr_block = GEN_3;
  assign io_out_bits_payload_client_xact_id = GEN_4;
  assign io_out_bits_payload_addr_beat = GEN_5;
  assign io_out_bits_payload_is_builtin_type = GEN_6;
  assign io_out_bits_payload_a_type = GEN_7;
  assign io_out_bits_payload_union = GEN_8;
  assign io_out_bits_payload_data = GEN_9;
  assign io_chosen = GEN_42;
  assign choice = GEN_49;
  assign GEN_0 = GEN_12;
  assign GEN_10 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_11 = 2'h2 == io_chosen ? io_in_2_valid : GEN_10;
  assign GEN_12 = 2'h3 == io_chosen ? io_in_3_valid : GEN_11;
  assign GEN_1 = GEN_15;
  assign GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_14 = 2'h2 == io_chosen ? io_in_2_bits_header_src : GEN_13;
  assign GEN_15 = 2'h3 == io_chosen ? io_in_3_bits_header_src : GEN_14;
  assign GEN_2 = GEN_18;
  assign GEN_16 = 2'h1 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_17 = 2'h2 == io_chosen ? io_in_2_bits_header_dst : GEN_16;
  assign GEN_18 = 2'h3 == io_chosen ? io_in_3_bits_header_dst : GEN_17;
  assign GEN_3 = GEN_21;
  assign GEN_19 = 2'h1 == io_chosen ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign GEN_20 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_block : GEN_19;
  assign GEN_21 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_block : GEN_20;
  assign GEN_4 = GEN_24;
  assign GEN_22 = 2'h1 == io_chosen ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign GEN_23 = 2'h2 == io_chosen ? io_in_2_bits_payload_client_xact_id : GEN_22;
  assign GEN_24 = 2'h3 == io_chosen ? io_in_3_bits_payload_client_xact_id : GEN_23;
  assign GEN_5 = GEN_27;
  assign GEN_25 = 2'h1 == io_chosen ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign GEN_26 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_beat : GEN_25;
  assign GEN_27 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_beat : GEN_26;
  assign GEN_6 = GEN_30;
  assign GEN_28 = 2'h1 == io_chosen ? io_in_1_bits_payload_is_builtin_type : io_in_0_bits_payload_is_builtin_type;
  assign GEN_29 = 2'h2 == io_chosen ? io_in_2_bits_payload_is_builtin_type : GEN_28;
  assign GEN_30 = 2'h3 == io_chosen ? io_in_3_bits_payload_is_builtin_type : GEN_29;
  assign GEN_7 = GEN_33;
  assign GEN_31 = 2'h1 == io_chosen ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign GEN_32 = 2'h2 == io_chosen ? io_in_2_bits_payload_a_type : GEN_31;
  assign GEN_33 = 2'h3 == io_chosen ? io_in_3_bits_payload_a_type : GEN_32;
  assign GEN_8 = GEN_36;
  assign GEN_34 = 2'h1 == io_chosen ? io_in_1_bits_payload_union : io_in_0_bits_payload_union;
  assign GEN_35 = 2'h2 == io_chosen ? io_in_2_bits_payload_union : GEN_34;
  assign GEN_36 = 2'h3 == io_chosen ? io_in_3_bits_payload_union : GEN_35;
  assign GEN_9 = GEN_39;
  assign GEN_37 = 2'h1 == io_chosen ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign GEN_38 = 2'h2 == io_chosen ? io_in_2_bits_payload_data : GEN_37;
  assign GEN_39 = 2'h3 == io_chosen ? io_in_3_bits_payload_data : GEN_38;
  assign T_1138 = T_1134 != 3'h0;
  assign T_1147_0 = 3'h3;
  assign T_1149 = io_out_bits_payload_a_type == T_1147_0;
  assign T_1150 = io_out_bits_payload_is_builtin_type & T_1149;
  assign T_1151 = io_out_ready & io_out_valid;
  assign T_1152 = T_1151 & T_1150;
  assign T_1156 = T_1134 + 3'h1;
  assign T_1157 = T_1156[2:0];
  assign GEN_40 = T_1152 ? io_chosen : T_1136;
  assign GEN_41 = T_1152 ? T_1157 : T_1134;
  assign GEN_42 = T_1138 ? T_1136 : choice;
  assign GEN_43 = T_1151 ? io_chosen : lastGrant;
  assign T_1162 = 2'h1 > lastGrant;
  assign T_1164 = 2'h2 > lastGrant;
  assign T_1166 = 2'h3 > lastGrant;
  assign T_1168 = io_in_1_valid & T_1162;
  assign T_1169 = io_in_2_valid & T_1164;
  assign T_1170 = io_in_3_valid & T_1166;
  assign T_1173 = T_1168 | T_1169;
  assign T_1174 = T_1173 | T_1170;
  assign T_1175 = T_1174 | io_in_0_valid;
  assign T_1176 = T_1175 | io_in_1_valid;
  assign T_1177 = T_1176 | io_in_2_valid;
  assign T_1181 = T_1168 == 1'h0;
  assign T_1183 = T_1173 == 1'h0;
  assign T_1185 = T_1174 == 1'h0;
  assign T_1187 = T_1175 == 1'h0;
  assign T_1189 = T_1176 == 1'h0;
  assign T_1191 = T_1177 == 1'h0;
  assign T_1195 = T_1162 | T_1187;
  assign T_1196 = T_1181 & T_1164;
  assign T_1197 = T_1196 | T_1189;
  assign T_1198 = T_1183 & T_1166;
  assign T_1199 = T_1198 | T_1191;
  assign T_1201 = T_1136 == 2'h0;
  assign T_1202 = T_1138 ? T_1201 : T_1185;
  assign T_1203 = T_1202 & io_out_ready;
  assign T_1205 = T_1136 == 2'h1;
  assign T_1206 = T_1138 ? T_1205 : T_1195;
  assign T_1207 = T_1206 & io_out_ready;
  assign T_1209 = T_1136 == 2'h2;
  assign T_1210 = T_1138 ? T_1209 : T_1197;
  assign T_1211 = T_1210 & io_out_ready;
  assign T_1213 = T_1136 == 2'h3;
  assign T_1214 = T_1138 ? T_1213 : T_1199;
  assign T_1215 = T_1214 & io_out_ready;
  assign GEN_44 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_45 = io_in_1_valid ? 2'h1 : GEN_44;
  assign GEN_46 = io_in_0_valid ? 2'h0 : GEN_45;
  assign GEN_47 = T_1170 ? 2'h3 : GEN_46;
  assign GEN_48 = T_1169 ? 2'h2 : GEN_47;
  assign GEN_49 = T_1168 ? 2'h1 : GEN_48;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_50 = {1{$random}};
  T_1134 = GEN_50[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_51 = {1{$random}};
  T_1136 = GEN_51[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_52 = {1{$random}};
  lastGrant = GEN_52[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1134 <= 3'h0;
    end else begin
      if(T_1152) begin
        T_1134 <= T_1157;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1152) begin
        T_1136 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1151) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module BasicBus(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input   io_in_0_bits_payload_client_xact_id,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input   io_in_0_bits_payload_is_builtin_type,
  input  [2:0] io_in_0_bits_payload_a_type,
  input  [11:0] io_in_0_bits_payload_union,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input   io_in_1_bits_payload_client_xact_id,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input   io_in_1_bits_payload_is_builtin_type,
  input  [2:0] io_in_1_bits_payload_a_type,
  input  [11:0] io_in_1_bits_payload_union,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input   io_in_2_bits_payload_client_xact_id,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input   io_in_2_bits_payload_is_builtin_type,
  input  [2:0] io_in_2_bits_payload_a_type,
  input  [11:0] io_in_2_bits_payload_union,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input   io_in_3_bits_payload_client_xact_id,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input   io_in_3_bits_payload_is_builtin_type,
  input  [2:0] io_in_3_bits_payload_a_type,
  input  [11:0] io_in_3_bits_payload_union,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [1:0] io_out_0_bits_header_src,
  output [1:0] io_out_0_bits_header_dst,
  output [25:0] io_out_0_bits_payload_addr_block,
  output  io_out_0_bits_payload_client_xact_id,
  output [2:0] io_out_0_bits_payload_addr_beat,
  output  io_out_0_bits_payload_is_builtin_type,
  output [2:0] io_out_0_bits_payload_a_type,
  output [11:0] io_out_0_bits_payload_union,
  output [63:0] io_out_0_bits_payload_data,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [1:0] io_out_1_bits_header_src,
  output [1:0] io_out_1_bits_header_dst,
  output [25:0] io_out_1_bits_payload_addr_block,
  output  io_out_1_bits_payload_client_xact_id,
  output [2:0] io_out_1_bits_payload_addr_beat,
  output  io_out_1_bits_payload_is_builtin_type,
  output [2:0] io_out_1_bits_payload_a_type,
  output [11:0] io_out_1_bits_payload_union,
  output [63:0] io_out_1_bits_payload_data,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [1:0] io_out_2_bits_header_src,
  output [1:0] io_out_2_bits_header_dst,
  output [25:0] io_out_2_bits_payload_addr_block,
  output  io_out_2_bits_payload_client_xact_id,
  output [2:0] io_out_2_bits_payload_addr_beat,
  output  io_out_2_bits_payload_is_builtin_type,
  output [2:0] io_out_2_bits_payload_a_type,
  output [11:0] io_out_2_bits_payload_union,
  output [63:0] io_out_2_bits_payload_data,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [1:0] io_out_3_bits_header_src,
  output [1:0] io_out_3_bits_header_dst,
  output [25:0] io_out_3_bits_payload_addr_block,
  output  io_out_3_bits_payload_client_xact_id,
  output [2:0] io_out_3_bits_payload_addr_beat,
  output  io_out_3_bits_payload_is_builtin_type,
  output [2:0] io_out_3_bits_payload_a_type,
  output [11:0] io_out_3_bits_payload_union,
  output [63:0] io_out_3_bits_payload_data
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_header_src;
  wire [1:0] arb_io_in_0_bits_header_dst;
  wire [25:0] arb_io_in_0_bits_payload_addr_block;
  wire  arb_io_in_0_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_0_bits_payload_addr_beat;
  wire  arb_io_in_0_bits_payload_is_builtin_type;
  wire [2:0] arb_io_in_0_bits_payload_a_type;
  wire [11:0] arb_io_in_0_bits_payload_union;
  wire [63:0] arb_io_in_0_bits_payload_data;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_header_src;
  wire [1:0] arb_io_in_1_bits_header_dst;
  wire [25:0] arb_io_in_1_bits_payload_addr_block;
  wire  arb_io_in_1_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_1_bits_payload_addr_beat;
  wire  arb_io_in_1_bits_payload_is_builtin_type;
  wire [2:0] arb_io_in_1_bits_payload_a_type;
  wire [11:0] arb_io_in_1_bits_payload_union;
  wire [63:0] arb_io_in_1_bits_payload_data;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [1:0] arb_io_in_2_bits_header_src;
  wire [1:0] arb_io_in_2_bits_header_dst;
  wire [25:0] arb_io_in_2_bits_payload_addr_block;
  wire  arb_io_in_2_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_2_bits_payload_addr_beat;
  wire  arb_io_in_2_bits_payload_is_builtin_type;
  wire [2:0] arb_io_in_2_bits_payload_a_type;
  wire [11:0] arb_io_in_2_bits_payload_union;
  wire [63:0] arb_io_in_2_bits_payload_data;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [1:0] arb_io_in_3_bits_header_src;
  wire [1:0] arb_io_in_3_bits_header_dst;
  wire [25:0] arb_io_in_3_bits_payload_addr_block;
  wire  arb_io_in_3_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_3_bits_payload_addr_beat;
  wire  arb_io_in_3_bits_payload_is_builtin_type;
  wire [2:0] arb_io_in_3_bits_payload_a_type;
  wire [11:0] arb_io_in_3_bits_payload_union;
  wire [63:0] arb_io_in_3_bits_payload_data;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_header_src;
  wire [1:0] arb_io_out_bits_header_dst;
  wire [25:0] arb_io_out_bits_payload_addr_block;
  wire  arb_io_out_bits_payload_client_xact_id;
  wire [2:0] arb_io_out_bits_payload_addr_beat;
  wire  arb_io_out_bits_payload_is_builtin_type;
  wire [2:0] arb_io_out_bits_payload_a_type;
  wire [11:0] arb_io_out_bits_payload_union;
  wire [63:0] arb_io_out_bits_payload_data;
  wire [1:0] arb_io_chosen;
  wire  GEN_0;
  wire  GEN_1;
  wire  GEN_2;
  wire  GEN_3;
  wire  T_1529;
  wire  T_1530;
  wire  T_1532;
  wire  T_1533;
  wire  T_1535;
  wire  T_1536;
  wire  T_1538;
  wire  T_1539;
  LockingRRArbiter arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_block(arb_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_client_xact_id(arb_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_addr_beat(arb_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_is_builtin_type(arb_io_in_0_bits_payload_is_builtin_type),
    .io_in_0_bits_payload_a_type(arb_io_in_0_bits_payload_a_type),
    .io_in_0_bits_payload_union(arb_io_in_0_bits_payload_union),
    .io_in_0_bits_payload_data(arb_io_in_0_bits_payload_data),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_block(arb_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_client_xact_id(arb_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_addr_beat(arb_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_is_builtin_type(arb_io_in_1_bits_payload_is_builtin_type),
    .io_in_1_bits_payload_a_type(arb_io_in_1_bits_payload_a_type),
    .io_in_1_bits_payload_union(arb_io_in_1_bits_payload_union),
    .io_in_1_bits_payload_data(arb_io_in_1_bits_payload_data),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_block(arb_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_client_xact_id(arb_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_addr_beat(arb_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_is_builtin_type(arb_io_in_2_bits_payload_is_builtin_type),
    .io_in_2_bits_payload_a_type(arb_io_in_2_bits_payload_a_type),
    .io_in_2_bits_payload_union(arb_io_in_2_bits_payload_union),
    .io_in_2_bits_payload_data(arb_io_in_2_bits_payload_data),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_block(arb_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_client_xact_id(arb_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_addr_beat(arb_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_is_builtin_type(arb_io_in_3_bits_payload_is_builtin_type),
    .io_in_3_bits_payload_a_type(arb_io_in_3_bits_payload_a_type),
    .io_in_3_bits_payload_union(arb_io_in_3_bits_payload_union),
    .io_in_3_bits_payload_data(arb_io_in_3_bits_payload_data),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_addr_block(arb_io_out_bits_payload_addr_block),
    .io_out_bits_payload_client_xact_id(arb_io_out_bits_payload_client_xact_id),
    .io_out_bits_payload_addr_beat(arb_io_out_bits_payload_addr_beat),
    .io_out_bits_payload_is_builtin_type(arb_io_out_bits_payload_is_builtin_type),
    .io_out_bits_payload_a_type(arb_io_out_bits_payload_a_type),
    .io_out_bits_payload_union(arb_io_out_bits_payload_union),
    .io_out_bits_payload_data(arb_io_out_bits_payload_data),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_out_0_valid = T_1530;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_0_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_0_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_0_bits_payload_a_type = arb_io_out_bits_payload_a_type;
  assign io_out_0_bits_payload_union = arb_io_out_bits_payload_union;
  assign io_out_0_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_1_valid = T_1533;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_1_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_1_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_1_bits_payload_a_type = arb_io_out_bits_payload_a_type;
  assign io_out_1_bits_payload_union = arb_io_out_bits_payload_union;
  assign io_out_1_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_2_valid = T_1536;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_2_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_2_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_2_bits_payload_a_type = arb_io_out_bits_payload_a_type;
  assign io_out_2_bits_payload_union = arb_io_out_bits_payload_union;
  assign io_out_2_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_3_valid = T_1539;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_3_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_3_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_3_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_3_bits_payload_a_type = arb_io_out_bits_payload_a_type;
  assign io_out_3_bits_payload_union = arb_io_out_bits_payload_union;
  assign io_out_3_bits_payload_data = arb_io_out_bits_payload_data;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_addr_block = io_in_0_bits_payload_addr_block;
  assign arb_io_in_0_bits_payload_client_xact_id = io_in_0_bits_payload_client_xact_id;
  assign arb_io_in_0_bits_payload_addr_beat = io_in_0_bits_payload_addr_beat;
  assign arb_io_in_0_bits_payload_is_builtin_type = io_in_0_bits_payload_is_builtin_type;
  assign arb_io_in_0_bits_payload_a_type = io_in_0_bits_payload_a_type;
  assign arb_io_in_0_bits_payload_union = io_in_0_bits_payload_union;
  assign arb_io_in_0_bits_payload_data = io_in_0_bits_payload_data;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_addr_block = io_in_1_bits_payload_addr_block;
  assign arb_io_in_1_bits_payload_client_xact_id = io_in_1_bits_payload_client_xact_id;
  assign arb_io_in_1_bits_payload_addr_beat = io_in_1_bits_payload_addr_beat;
  assign arb_io_in_1_bits_payload_is_builtin_type = io_in_1_bits_payload_is_builtin_type;
  assign arb_io_in_1_bits_payload_a_type = io_in_1_bits_payload_a_type;
  assign arb_io_in_1_bits_payload_union = io_in_1_bits_payload_union;
  assign arb_io_in_1_bits_payload_data = io_in_1_bits_payload_data;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_addr_block = io_in_2_bits_payload_addr_block;
  assign arb_io_in_2_bits_payload_client_xact_id = io_in_2_bits_payload_client_xact_id;
  assign arb_io_in_2_bits_payload_addr_beat = io_in_2_bits_payload_addr_beat;
  assign arb_io_in_2_bits_payload_is_builtin_type = io_in_2_bits_payload_is_builtin_type;
  assign arb_io_in_2_bits_payload_a_type = io_in_2_bits_payload_a_type;
  assign arb_io_in_2_bits_payload_union = io_in_2_bits_payload_union;
  assign arb_io_in_2_bits_payload_data = io_in_2_bits_payload_data;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_addr_block = io_in_3_bits_payload_addr_block;
  assign arb_io_in_3_bits_payload_client_xact_id = io_in_3_bits_payload_client_xact_id;
  assign arb_io_in_3_bits_payload_addr_beat = io_in_3_bits_payload_addr_beat;
  assign arb_io_in_3_bits_payload_is_builtin_type = io_in_3_bits_payload_is_builtin_type;
  assign arb_io_in_3_bits_payload_a_type = io_in_3_bits_payload_a_type;
  assign arb_io_in_3_bits_payload_union = io_in_3_bits_payload_union;
  assign arb_io_in_3_bits_payload_data = io_in_3_bits_payload_data;
  assign arb_io_out_ready = GEN_0;
  assign GEN_0 = GEN_3;
  assign GEN_1 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_2 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_3 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_2;
  assign T_1529 = arb_io_out_bits_header_dst == 2'h0;
  assign T_1530 = arb_io_out_valid & T_1529;
  assign T_1532 = arb_io_out_bits_header_dst == 2'h1;
  assign T_1533 = arb_io_out_valid & T_1532;
  assign T_1535 = arb_io_out_bits_header_dst == 2'h2;
  assign T_1536 = arb_io_out_valid & T_1535;
  assign T_1538 = arb_io_out_bits_header_dst == 2'h3;
  assign T_1539 = arb_io_out_valid & T_1538;
endmodule
module LockingRRArbiter_1(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input   io_in_0_bits_payload_client_xact_id,
  input   io_in_0_bits_payload_voluntary,
  input  [2:0] io_in_0_bits_payload_r_type,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input   io_in_1_bits_payload_client_xact_id,
  input   io_in_1_bits_payload_voluntary,
  input  [2:0] io_in_1_bits_payload_r_type,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input   io_in_2_bits_payload_client_xact_id,
  input   io_in_2_bits_payload_voluntary,
  input  [2:0] io_in_2_bits_payload_r_type,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input   io_in_3_bits_payload_client_xact_id,
  input   io_in_3_bits_payload_voluntary,
  input  [2:0] io_in_3_bits_payload_r_type,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_ready,
  output  io_out_valid,
  output [1:0] io_out_bits_header_src,
  output [1:0] io_out_bits_header_dst,
  output [2:0] io_out_bits_payload_addr_beat,
  output [25:0] io_out_bits_payload_addr_block,
  output  io_out_bits_payload_client_xact_id,
  output  io_out_bits_payload_voluntary,
  output [2:0] io_out_bits_payload_r_type,
  output [63:0] io_out_bits_payload_data,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire [1:0] GEN_1;
  wire [1:0] GEN_12;
  wire [1:0] GEN_13;
  wire [1:0] GEN_14;
  wire [1:0] GEN_2;
  wire [1:0] GEN_15;
  wire [1:0] GEN_16;
  wire [1:0] GEN_17;
  wire [2:0] GEN_3;
  wire [2:0] GEN_18;
  wire [2:0] GEN_19;
  wire [2:0] GEN_20;
  wire [25:0] GEN_4;
  wire [25:0] GEN_21;
  wire [25:0] GEN_22;
  wire [25:0] GEN_23;
  wire  GEN_5;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_6;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_29;
  wire [2:0] GEN_7;
  wire [2:0] GEN_30;
  wire [2:0] GEN_31;
  wire [2:0] GEN_32;
  wire [63:0] GEN_8;
  wire [63:0] GEN_33;
  wire [63:0] GEN_34;
  wire [63:0] GEN_35;
  reg [2:0] T_1100;
  reg [31:0] GEN_46;
  reg [1:0] T_1102;
  reg [31:0] GEN_47;
  wire  T_1104;
  wire  T_1106;
  wire  T_1107;
  wire  T_1108;
  wire  T_1109;
  wire  T_1110;
  wire  T_1112;
  wire  T_1113;
  wire [3:0] T_1117;
  wire [2:0] T_1118;
  wire [1:0] GEN_36;
  wire [2:0] GEN_37;
  wire [1:0] GEN_38;
  reg [1:0] lastGrant;
  reg [31:0] GEN_48;
  wire [1:0] GEN_39;
  wire  T_1123;
  wire  T_1125;
  wire  T_1127;
  wire  T_1129;
  wire  T_1130;
  wire  T_1131;
  wire  T_1134;
  wire  T_1135;
  wire  T_1136;
  wire  T_1137;
  wire  T_1138;
  wire  T_1142;
  wire  T_1144;
  wire  T_1146;
  wire  T_1148;
  wire  T_1150;
  wire  T_1152;
  wire  T_1156;
  wire  T_1157;
  wire  T_1158;
  wire  T_1159;
  wire  T_1160;
  wire  T_1162;
  wire  T_1163;
  wire  T_1164;
  wire  T_1166;
  wire  T_1167;
  wire  T_1168;
  wire  T_1170;
  wire  T_1171;
  wire  T_1172;
  wire  T_1174;
  wire  T_1175;
  wire  T_1176;
  wire [1:0] GEN_40;
  wire [1:0] GEN_41;
  wire [1:0] GEN_42;
  wire [1:0] GEN_43;
  wire [1:0] GEN_44;
  wire [1:0] GEN_45;
  assign io_in_0_ready = T_1164;
  assign io_in_1_ready = T_1168;
  assign io_in_2_ready = T_1172;
  assign io_in_3_ready = T_1176;
  assign io_out_valid = GEN_0;
  assign io_out_bits_header_src = GEN_1;
  assign io_out_bits_header_dst = GEN_2;
  assign io_out_bits_payload_addr_beat = GEN_3;
  assign io_out_bits_payload_addr_block = GEN_4;
  assign io_out_bits_payload_client_xact_id = GEN_5;
  assign io_out_bits_payload_voluntary = GEN_6;
  assign io_out_bits_payload_r_type = GEN_7;
  assign io_out_bits_payload_data = GEN_8;
  assign io_chosen = GEN_38;
  assign choice = GEN_45;
  assign GEN_0 = GEN_11;
  assign GEN_9 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_10 = 2'h2 == io_chosen ? io_in_2_valid : GEN_9;
  assign GEN_11 = 2'h3 == io_chosen ? io_in_3_valid : GEN_10;
  assign GEN_1 = GEN_14;
  assign GEN_12 = 2'h1 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_13 = 2'h2 == io_chosen ? io_in_2_bits_header_src : GEN_12;
  assign GEN_14 = 2'h3 == io_chosen ? io_in_3_bits_header_src : GEN_13;
  assign GEN_2 = GEN_17;
  assign GEN_15 = 2'h1 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_16 = 2'h2 == io_chosen ? io_in_2_bits_header_dst : GEN_15;
  assign GEN_17 = 2'h3 == io_chosen ? io_in_3_bits_header_dst : GEN_16;
  assign GEN_3 = GEN_20;
  assign GEN_18 = 2'h1 == io_chosen ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign GEN_19 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_beat : GEN_18;
  assign GEN_20 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_beat : GEN_19;
  assign GEN_4 = GEN_23;
  assign GEN_21 = 2'h1 == io_chosen ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_block : GEN_21;
  assign GEN_23 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_block : GEN_22;
  assign GEN_5 = GEN_26;
  assign GEN_24 = 2'h1 == io_chosen ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign GEN_25 = 2'h2 == io_chosen ? io_in_2_bits_payload_client_xact_id : GEN_24;
  assign GEN_26 = 2'h3 == io_chosen ? io_in_3_bits_payload_client_xact_id : GEN_25;
  assign GEN_6 = GEN_29;
  assign GEN_27 = 2'h1 == io_chosen ? io_in_1_bits_payload_voluntary : io_in_0_bits_payload_voluntary;
  assign GEN_28 = 2'h2 == io_chosen ? io_in_2_bits_payload_voluntary : GEN_27;
  assign GEN_29 = 2'h3 == io_chosen ? io_in_3_bits_payload_voluntary : GEN_28;
  assign GEN_7 = GEN_32;
  assign GEN_30 = 2'h1 == io_chosen ? io_in_1_bits_payload_r_type : io_in_0_bits_payload_r_type;
  assign GEN_31 = 2'h2 == io_chosen ? io_in_2_bits_payload_r_type : GEN_30;
  assign GEN_32 = 2'h3 == io_chosen ? io_in_3_bits_payload_r_type : GEN_31;
  assign GEN_8 = GEN_35;
  assign GEN_33 = 2'h1 == io_chosen ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign GEN_34 = 2'h2 == io_chosen ? io_in_2_bits_payload_data : GEN_33;
  assign GEN_35 = 2'h3 == io_chosen ? io_in_3_bits_payload_data : GEN_34;
  assign T_1104 = T_1100 != 3'h0;
  assign T_1106 = io_out_bits_payload_r_type == 3'h0;
  assign T_1107 = io_out_bits_payload_r_type == 3'h1;
  assign T_1108 = io_out_bits_payload_r_type == 3'h2;
  assign T_1109 = T_1106 | T_1107;
  assign T_1110 = T_1109 | T_1108;
  assign T_1112 = io_out_ready & io_out_valid;
  assign T_1113 = T_1112 & T_1110;
  assign T_1117 = T_1100 + 3'h1;
  assign T_1118 = T_1117[2:0];
  assign GEN_36 = T_1113 ? io_chosen : T_1102;
  assign GEN_37 = T_1113 ? T_1118 : T_1100;
  assign GEN_38 = T_1104 ? T_1102 : choice;
  assign GEN_39 = T_1112 ? io_chosen : lastGrant;
  assign T_1123 = 2'h1 > lastGrant;
  assign T_1125 = 2'h2 > lastGrant;
  assign T_1127 = 2'h3 > lastGrant;
  assign T_1129 = io_in_1_valid & T_1123;
  assign T_1130 = io_in_2_valid & T_1125;
  assign T_1131 = io_in_3_valid & T_1127;
  assign T_1134 = T_1129 | T_1130;
  assign T_1135 = T_1134 | T_1131;
  assign T_1136 = T_1135 | io_in_0_valid;
  assign T_1137 = T_1136 | io_in_1_valid;
  assign T_1138 = T_1137 | io_in_2_valid;
  assign T_1142 = T_1129 == 1'h0;
  assign T_1144 = T_1134 == 1'h0;
  assign T_1146 = T_1135 == 1'h0;
  assign T_1148 = T_1136 == 1'h0;
  assign T_1150 = T_1137 == 1'h0;
  assign T_1152 = T_1138 == 1'h0;
  assign T_1156 = T_1123 | T_1148;
  assign T_1157 = T_1142 & T_1125;
  assign T_1158 = T_1157 | T_1150;
  assign T_1159 = T_1144 & T_1127;
  assign T_1160 = T_1159 | T_1152;
  assign T_1162 = T_1102 == 2'h0;
  assign T_1163 = T_1104 ? T_1162 : T_1146;
  assign T_1164 = T_1163 & io_out_ready;
  assign T_1166 = T_1102 == 2'h1;
  assign T_1167 = T_1104 ? T_1166 : T_1156;
  assign T_1168 = T_1167 & io_out_ready;
  assign T_1170 = T_1102 == 2'h2;
  assign T_1171 = T_1104 ? T_1170 : T_1158;
  assign T_1172 = T_1171 & io_out_ready;
  assign T_1174 = T_1102 == 2'h3;
  assign T_1175 = T_1104 ? T_1174 : T_1160;
  assign T_1176 = T_1175 & io_out_ready;
  assign GEN_40 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_41 = io_in_1_valid ? 2'h1 : GEN_40;
  assign GEN_42 = io_in_0_valid ? 2'h0 : GEN_41;
  assign GEN_43 = T_1131 ? 2'h3 : GEN_42;
  assign GEN_44 = T_1130 ? 2'h2 : GEN_43;
  assign GEN_45 = T_1129 ? 2'h1 : GEN_44;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_46 = {1{$random}};
  T_1100 = GEN_46[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_47 = {1{$random}};
  T_1102 = GEN_47[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_48 = {1{$random}};
  lastGrant = GEN_48[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1100 <= 3'h0;
    end else begin
      if(T_1113) begin
        T_1100 <= T_1118;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1113) begin
        T_1102 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1112) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module BasicBus_1(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input   io_in_0_bits_payload_client_xact_id,
  input   io_in_0_bits_payload_voluntary,
  input  [2:0] io_in_0_bits_payload_r_type,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input   io_in_1_bits_payload_client_xact_id,
  input   io_in_1_bits_payload_voluntary,
  input  [2:0] io_in_1_bits_payload_r_type,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input   io_in_2_bits_payload_client_xact_id,
  input   io_in_2_bits_payload_voluntary,
  input  [2:0] io_in_2_bits_payload_r_type,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input   io_in_3_bits_payload_client_xact_id,
  input   io_in_3_bits_payload_voluntary,
  input  [2:0] io_in_3_bits_payload_r_type,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [1:0] io_out_0_bits_header_src,
  output [1:0] io_out_0_bits_header_dst,
  output [2:0] io_out_0_bits_payload_addr_beat,
  output [25:0] io_out_0_bits_payload_addr_block,
  output  io_out_0_bits_payload_client_xact_id,
  output  io_out_0_bits_payload_voluntary,
  output [2:0] io_out_0_bits_payload_r_type,
  output [63:0] io_out_0_bits_payload_data,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [1:0] io_out_1_bits_header_src,
  output [1:0] io_out_1_bits_header_dst,
  output [2:0] io_out_1_bits_payload_addr_beat,
  output [25:0] io_out_1_bits_payload_addr_block,
  output  io_out_1_bits_payload_client_xact_id,
  output  io_out_1_bits_payload_voluntary,
  output [2:0] io_out_1_bits_payload_r_type,
  output [63:0] io_out_1_bits_payload_data,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [1:0] io_out_2_bits_header_src,
  output [1:0] io_out_2_bits_header_dst,
  output [2:0] io_out_2_bits_payload_addr_beat,
  output [25:0] io_out_2_bits_payload_addr_block,
  output  io_out_2_bits_payload_client_xact_id,
  output  io_out_2_bits_payload_voluntary,
  output [2:0] io_out_2_bits_payload_r_type,
  output [63:0] io_out_2_bits_payload_data,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [1:0] io_out_3_bits_header_src,
  output [1:0] io_out_3_bits_header_dst,
  output [2:0] io_out_3_bits_payload_addr_beat,
  output [25:0] io_out_3_bits_payload_addr_block,
  output  io_out_3_bits_payload_client_xact_id,
  output  io_out_3_bits_payload_voluntary,
  output [2:0] io_out_3_bits_payload_r_type,
  output [63:0] io_out_3_bits_payload_data
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_header_src;
  wire [1:0] arb_io_in_0_bits_header_dst;
  wire [2:0] arb_io_in_0_bits_payload_addr_beat;
  wire [25:0] arb_io_in_0_bits_payload_addr_block;
  wire  arb_io_in_0_bits_payload_client_xact_id;
  wire  arb_io_in_0_bits_payload_voluntary;
  wire [2:0] arb_io_in_0_bits_payload_r_type;
  wire [63:0] arb_io_in_0_bits_payload_data;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_header_src;
  wire [1:0] arb_io_in_1_bits_header_dst;
  wire [2:0] arb_io_in_1_bits_payload_addr_beat;
  wire [25:0] arb_io_in_1_bits_payload_addr_block;
  wire  arb_io_in_1_bits_payload_client_xact_id;
  wire  arb_io_in_1_bits_payload_voluntary;
  wire [2:0] arb_io_in_1_bits_payload_r_type;
  wire [63:0] arb_io_in_1_bits_payload_data;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [1:0] arb_io_in_2_bits_header_src;
  wire [1:0] arb_io_in_2_bits_header_dst;
  wire [2:0] arb_io_in_2_bits_payload_addr_beat;
  wire [25:0] arb_io_in_2_bits_payload_addr_block;
  wire  arb_io_in_2_bits_payload_client_xact_id;
  wire  arb_io_in_2_bits_payload_voluntary;
  wire [2:0] arb_io_in_2_bits_payload_r_type;
  wire [63:0] arb_io_in_2_bits_payload_data;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [1:0] arb_io_in_3_bits_header_src;
  wire [1:0] arb_io_in_3_bits_header_dst;
  wire [2:0] arb_io_in_3_bits_payload_addr_beat;
  wire [25:0] arb_io_in_3_bits_payload_addr_block;
  wire  arb_io_in_3_bits_payload_client_xact_id;
  wire  arb_io_in_3_bits_payload_voluntary;
  wire [2:0] arb_io_in_3_bits_payload_r_type;
  wire [63:0] arb_io_in_3_bits_payload_data;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_header_src;
  wire [1:0] arb_io_out_bits_header_dst;
  wire [2:0] arb_io_out_bits_payload_addr_beat;
  wire [25:0] arb_io_out_bits_payload_addr_block;
  wire  arb_io_out_bits_payload_client_xact_id;
  wire  arb_io_out_bits_payload_voluntary;
  wire [2:0] arb_io_out_bits_payload_r_type;
  wire [63:0] arb_io_out_bits_payload_data;
  wire [1:0] arb_io_chosen;
  wire  GEN_0;
  wire  GEN_1;
  wire  GEN_2;
  wire  GEN_3;
  wire  T_1483;
  wire  T_1484;
  wire  T_1486;
  wire  T_1487;
  wire  T_1489;
  wire  T_1490;
  wire  T_1492;
  wire  T_1493;
  LockingRRArbiter_1 arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_beat(arb_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_addr_block(arb_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_client_xact_id(arb_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_voluntary(arb_io_in_0_bits_payload_voluntary),
    .io_in_0_bits_payload_r_type(arb_io_in_0_bits_payload_r_type),
    .io_in_0_bits_payload_data(arb_io_in_0_bits_payload_data),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_beat(arb_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_addr_block(arb_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_client_xact_id(arb_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_voluntary(arb_io_in_1_bits_payload_voluntary),
    .io_in_1_bits_payload_r_type(arb_io_in_1_bits_payload_r_type),
    .io_in_1_bits_payload_data(arb_io_in_1_bits_payload_data),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_beat(arb_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_addr_block(arb_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_client_xact_id(arb_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_voluntary(arb_io_in_2_bits_payload_voluntary),
    .io_in_2_bits_payload_r_type(arb_io_in_2_bits_payload_r_type),
    .io_in_2_bits_payload_data(arb_io_in_2_bits_payload_data),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_beat(arb_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_addr_block(arb_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_client_xact_id(arb_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_voluntary(arb_io_in_3_bits_payload_voluntary),
    .io_in_3_bits_payload_r_type(arb_io_in_3_bits_payload_r_type),
    .io_in_3_bits_payload_data(arb_io_in_3_bits_payload_data),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_addr_beat(arb_io_out_bits_payload_addr_beat),
    .io_out_bits_payload_addr_block(arb_io_out_bits_payload_addr_block),
    .io_out_bits_payload_client_xact_id(arb_io_out_bits_payload_client_xact_id),
    .io_out_bits_payload_voluntary(arb_io_out_bits_payload_voluntary),
    .io_out_bits_payload_r_type(arb_io_out_bits_payload_r_type),
    .io_out_bits_payload_data(arb_io_out_bits_payload_data),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_out_0_valid = T_1484;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_0_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_0_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_voluntary = arb_io_out_bits_payload_voluntary;
  assign io_out_0_bits_payload_r_type = arb_io_out_bits_payload_r_type;
  assign io_out_0_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_1_valid = T_1487;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_1_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_1_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_voluntary = arb_io_out_bits_payload_voluntary;
  assign io_out_1_bits_payload_r_type = arb_io_out_bits_payload_r_type;
  assign io_out_1_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_2_valid = T_1490;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_2_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_2_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_voluntary = arb_io_out_bits_payload_voluntary;
  assign io_out_2_bits_payload_r_type = arb_io_out_bits_payload_r_type;
  assign io_out_2_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_3_valid = T_1493;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_3_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_3_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_3_bits_payload_voluntary = arb_io_out_bits_payload_voluntary;
  assign io_out_3_bits_payload_r_type = arb_io_out_bits_payload_r_type;
  assign io_out_3_bits_payload_data = arb_io_out_bits_payload_data;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_addr_beat = io_in_0_bits_payload_addr_beat;
  assign arb_io_in_0_bits_payload_addr_block = io_in_0_bits_payload_addr_block;
  assign arb_io_in_0_bits_payload_client_xact_id = io_in_0_bits_payload_client_xact_id;
  assign arb_io_in_0_bits_payload_voluntary = io_in_0_bits_payload_voluntary;
  assign arb_io_in_0_bits_payload_r_type = io_in_0_bits_payload_r_type;
  assign arb_io_in_0_bits_payload_data = io_in_0_bits_payload_data;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_addr_beat = io_in_1_bits_payload_addr_beat;
  assign arb_io_in_1_bits_payload_addr_block = io_in_1_bits_payload_addr_block;
  assign arb_io_in_1_bits_payload_client_xact_id = io_in_1_bits_payload_client_xact_id;
  assign arb_io_in_1_bits_payload_voluntary = io_in_1_bits_payload_voluntary;
  assign arb_io_in_1_bits_payload_r_type = io_in_1_bits_payload_r_type;
  assign arb_io_in_1_bits_payload_data = io_in_1_bits_payload_data;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_addr_beat = io_in_2_bits_payload_addr_beat;
  assign arb_io_in_2_bits_payload_addr_block = io_in_2_bits_payload_addr_block;
  assign arb_io_in_2_bits_payload_client_xact_id = io_in_2_bits_payload_client_xact_id;
  assign arb_io_in_2_bits_payload_voluntary = io_in_2_bits_payload_voluntary;
  assign arb_io_in_2_bits_payload_r_type = io_in_2_bits_payload_r_type;
  assign arb_io_in_2_bits_payload_data = io_in_2_bits_payload_data;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_addr_beat = io_in_3_bits_payload_addr_beat;
  assign arb_io_in_3_bits_payload_addr_block = io_in_3_bits_payload_addr_block;
  assign arb_io_in_3_bits_payload_client_xact_id = io_in_3_bits_payload_client_xact_id;
  assign arb_io_in_3_bits_payload_voluntary = io_in_3_bits_payload_voluntary;
  assign arb_io_in_3_bits_payload_r_type = io_in_3_bits_payload_r_type;
  assign arb_io_in_3_bits_payload_data = io_in_3_bits_payload_data;
  assign arb_io_out_ready = GEN_0;
  assign GEN_0 = GEN_3;
  assign GEN_1 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_2 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_3 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_2;
  assign T_1483 = arb_io_out_bits_header_dst == 2'h0;
  assign T_1484 = arb_io_out_valid & T_1483;
  assign T_1486 = arb_io_out_bits_header_dst == 2'h1;
  assign T_1487 = arb_io_out_valid & T_1486;
  assign T_1489 = arb_io_out_bits_header_dst == 2'h2;
  assign T_1490 = arb_io_out_valid & T_1489;
  assign T_1492 = arb_io_out_bits_header_dst == 2'h3;
  assign T_1493 = arb_io_out_valid & T_1492;
endmodule
module LockingRRArbiter_2(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_p_type,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_p_type,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_p_type,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_p_type,
  input   io_out_ready,
  output  io_out_valid,
  output [1:0] io_out_bits_header_src,
  output [1:0] io_out_bits_header_dst,
  output [25:0] io_out_bits_payload_addr_block,
  output [1:0] io_out_bits_payload_p_type,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire [1:0] GEN_1;
  wire [1:0] GEN_8;
  wire [1:0] GEN_9;
  wire [1:0] GEN_10;
  wire [1:0] GEN_2;
  wire [1:0] GEN_11;
  wire [1:0] GEN_12;
  wire [1:0] GEN_13;
  wire [25:0] GEN_3;
  wire [25:0] GEN_14;
  wire [25:0] GEN_15;
  wire [25:0] GEN_16;
  wire [1:0] GEN_4;
  wire [1:0] GEN_17;
  wire [1:0] GEN_18;
  wire [1:0] GEN_19;
  wire  T_964;
  reg [1:0] lastGrant;
  reg [31:0] GEN_27;
  wire [1:0] GEN_20;
  wire  T_967;
  wire  T_969;
  wire  T_971;
  wire  T_973;
  wire  T_974;
  wire  T_975;
  wire  T_978;
  wire  T_979;
  wire  T_980;
  wire  T_981;
  wire  T_982;
  wire  T_986;
  wire  T_988;
  wire  T_990;
  wire  T_992;
  wire  T_994;
  wire  T_996;
  wire  T_1000;
  wire  T_1001;
  wire  T_1002;
  wire  T_1003;
  wire  T_1004;
  wire  T_1005;
  wire  T_1006;
  wire  T_1007;
  wire  T_1008;
  wire [1:0] GEN_21;
  wire [1:0] GEN_22;
  wire [1:0] GEN_23;
  wire [1:0] GEN_24;
  wire [1:0] GEN_25;
  wire [1:0] GEN_26;
  assign io_in_0_ready = T_1005;
  assign io_in_1_ready = T_1006;
  assign io_in_2_ready = T_1007;
  assign io_in_3_ready = T_1008;
  assign io_out_valid = GEN_0;
  assign io_out_bits_header_src = GEN_1;
  assign io_out_bits_header_dst = GEN_2;
  assign io_out_bits_payload_addr_block = GEN_3;
  assign io_out_bits_payload_p_type = GEN_4;
  assign io_chosen = choice;
  assign choice = GEN_26;
  assign GEN_0 = GEN_7;
  assign GEN_5 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_6 = 2'h2 == io_chosen ? io_in_2_valid : GEN_5;
  assign GEN_7 = 2'h3 == io_chosen ? io_in_3_valid : GEN_6;
  assign GEN_1 = GEN_10;
  assign GEN_8 = 2'h1 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_9 = 2'h2 == io_chosen ? io_in_2_bits_header_src : GEN_8;
  assign GEN_10 = 2'h3 == io_chosen ? io_in_3_bits_header_src : GEN_9;
  assign GEN_2 = GEN_13;
  assign GEN_11 = 2'h1 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_12 = 2'h2 == io_chosen ? io_in_2_bits_header_dst : GEN_11;
  assign GEN_13 = 2'h3 == io_chosen ? io_in_3_bits_header_dst : GEN_12;
  assign GEN_3 = GEN_16;
  assign GEN_14 = 2'h1 == io_chosen ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign GEN_15 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_block : GEN_14;
  assign GEN_16 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_block : GEN_15;
  assign GEN_4 = GEN_19;
  assign GEN_17 = 2'h1 == io_chosen ? io_in_1_bits_payload_p_type : io_in_0_bits_payload_p_type;
  assign GEN_18 = 2'h2 == io_chosen ? io_in_2_bits_payload_p_type : GEN_17;
  assign GEN_19 = 2'h3 == io_chosen ? io_in_3_bits_payload_p_type : GEN_18;
  assign T_964 = io_out_ready & io_out_valid;
  assign GEN_20 = T_964 ? io_chosen : lastGrant;
  assign T_967 = 2'h1 > lastGrant;
  assign T_969 = 2'h2 > lastGrant;
  assign T_971 = 2'h3 > lastGrant;
  assign T_973 = io_in_1_valid & T_967;
  assign T_974 = io_in_2_valid & T_969;
  assign T_975 = io_in_3_valid & T_971;
  assign T_978 = T_973 | T_974;
  assign T_979 = T_978 | T_975;
  assign T_980 = T_979 | io_in_0_valid;
  assign T_981 = T_980 | io_in_1_valid;
  assign T_982 = T_981 | io_in_2_valid;
  assign T_986 = T_973 == 1'h0;
  assign T_988 = T_978 == 1'h0;
  assign T_990 = T_979 == 1'h0;
  assign T_992 = T_980 == 1'h0;
  assign T_994 = T_981 == 1'h0;
  assign T_996 = T_982 == 1'h0;
  assign T_1000 = T_967 | T_992;
  assign T_1001 = T_986 & T_969;
  assign T_1002 = T_1001 | T_994;
  assign T_1003 = T_988 & T_971;
  assign T_1004 = T_1003 | T_996;
  assign T_1005 = T_990 & io_out_ready;
  assign T_1006 = T_1000 & io_out_ready;
  assign T_1007 = T_1002 & io_out_ready;
  assign T_1008 = T_1004 & io_out_ready;
  assign GEN_21 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_22 = io_in_1_valid ? 2'h1 : GEN_21;
  assign GEN_23 = io_in_0_valid ? 2'h0 : GEN_22;
  assign GEN_24 = T_975 ? 2'h3 : GEN_23;
  assign GEN_25 = T_974 ? 2'h2 : GEN_24;
  assign GEN_26 = T_973 ? 2'h1 : GEN_25;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_27 = {1{$random}};
  lastGrant = GEN_27[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_964) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module BasicBus_2(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_p_type,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_p_type,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_p_type,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_p_type,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [1:0] io_out_0_bits_header_src,
  output [1:0] io_out_0_bits_header_dst,
  output [25:0] io_out_0_bits_payload_addr_block,
  output [1:0] io_out_0_bits_payload_p_type,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [1:0] io_out_1_bits_header_src,
  output [1:0] io_out_1_bits_header_dst,
  output [25:0] io_out_1_bits_payload_addr_block,
  output [1:0] io_out_1_bits_payload_p_type,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [1:0] io_out_2_bits_header_src,
  output [1:0] io_out_2_bits_header_dst,
  output [25:0] io_out_2_bits_payload_addr_block,
  output [1:0] io_out_2_bits_payload_p_type,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [1:0] io_out_3_bits_header_src,
  output [1:0] io_out_3_bits_header_dst,
  output [25:0] io_out_3_bits_payload_addr_block,
  output [1:0] io_out_3_bits_payload_p_type
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_header_src;
  wire [1:0] arb_io_in_0_bits_header_dst;
  wire [25:0] arb_io_in_0_bits_payload_addr_block;
  wire [1:0] arb_io_in_0_bits_payload_p_type;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_header_src;
  wire [1:0] arb_io_in_1_bits_header_dst;
  wire [25:0] arb_io_in_1_bits_payload_addr_block;
  wire [1:0] arb_io_in_1_bits_payload_p_type;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [1:0] arb_io_in_2_bits_header_src;
  wire [1:0] arb_io_in_2_bits_header_dst;
  wire [25:0] arb_io_in_2_bits_payload_addr_block;
  wire [1:0] arb_io_in_2_bits_payload_p_type;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [1:0] arb_io_in_3_bits_header_src;
  wire [1:0] arb_io_in_3_bits_header_dst;
  wire [25:0] arb_io_in_3_bits_payload_addr_block;
  wire [1:0] arb_io_in_3_bits_payload_p_type;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_header_src;
  wire [1:0] arb_io_out_bits_header_dst;
  wire [25:0] arb_io_out_bits_payload_addr_block;
  wire [1:0] arb_io_out_bits_payload_p_type;
  wire [1:0] arb_io_chosen;
  wire  GEN_0;
  wire  GEN_1;
  wire  GEN_2;
  wire  GEN_3;
  wire  T_1299;
  wire  T_1300;
  wire  T_1302;
  wire  T_1303;
  wire  T_1305;
  wire  T_1306;
  wire  T_1308;
  wire  T_1309;
  LockingRRArbiter_2 arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_block(arb_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_p_type(arb_io_in_0_bits_payload_p_type),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_block(arb_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_p_type(arb_io_in_1_bits_payload_p_type),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_block(arb_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_p_type(arb_io_in_2_bits_payload_p_type),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_block(arb_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_p_type(arb_io_in_3_bits_payload_p_type),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_addr_block(arb_io_out_bits_payload_addr_block),
    .io_out_bits_payload_p_type(arb_io_out_bits_payload_p_type),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_out_0_valid = T_1300;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_0_bits_payload_p_type = arb_io_out_bits_payload_p_type;
  assign io_out_1_valid = T_1303;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_1_bits_payload_p_type = arb_io_out_bits_payload_p_type;
  assign io_out_2_valid = T_1306;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_2_bits_payload_p_type = arb_io_out_bits_payload_p_type;
  assign io_out_3_valid = T_1309;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_3_bits_payload_p_type = arb_io_out_bits_payload_p_type;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_addr_block = io_in_0_bits_payload_addr_block;
  assign arb_io_in_0_bits_payload_p_type = io_in_0_bits_payload_p_type;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_addr_block = io_in_1_bits_payload_addr_block;
  assign arb_io_in_1_bits_payload_p_type = io_in_1_bits_payload_p_type;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_addr_block = io_in_2_bits_payload_addr_block;
  assign arb_io_in_2_bits_payload_p_type = io_in_2_bits_payload_p_type;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_addr_block = io_in_3_bits_payload_addr_block;
  assign arb_io_in_3_bits_payload_p_type = io_in_3_bits_payload_p_type;
  assign arb_io_out_ready = GEN_0;
  assign GEN_0 = GEN_3;
  assign GEN_1 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_2 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_3 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_2;
  assign T_1299 = arb_io_out_bits_header_dst == 2'h0;
  assign T_1300 = arb_io_out_valid & T_1299;
  assign T_1302 = arb_io_out_bits_header_dst == 2'h1;
  assign T_1303 = arb_io_out_valid & T_1302;
  assign T_1305 = arb_io_out_bits_header_dst == 2'h2;
  assign T_1306 = arb_io_out_valid & T_1305;
  assign T_1308 = arb_io_out_bits_header_dst == 2'h3;
  assign T_1309 = arb_io_out_valid & T_1308;
endmodule
module LockingRRArbiter_3(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input   io_in_0_bits_payload_client_xact_id,
  input  [1:0] io_in_0_bits_payload_manager_xact_id,
  input   io_in_0_bits_payload_is_builtin_type,
  input  [3:0] io_in_0_bits_payload_g_type,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input   io_in_1_bits_payload_client_xact_id,
  input  [1:0] io_in_1_bits_payload_manager_xact_id,
  input   io_in_1_bits_payload_is_builtin_type,
  input  [3:0] io_in_1_bits_payload_g_type,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input   io_in_2_bits_payload_client_xact_id,
  input  [1:0] io_in_2_bits_payload_manager_xact_id,
  input   io_in_2_bits_payload_is_builtin_type,
  input  [3:0] io_in_2_bits_payload_g_type,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input   io_in_3_bits_payload_client_xact_id,
  input  [1:0] io_in_3_bits_payload_manager_xact_id,
  input   io_in_3_bits_payload_is_builtin_type,
  input  [3:0] io_in_3_bits_payload_g_type,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_ready,
  output  io_out_valid,
  output [1:0] io_out_bits_header_src,
  output [1:0] io_out_bits_header_dst,
  output [2:0] io_out_bits_payload_addr_beat,
  output  io_out_bits_payload_client_xact_id,
  output [1:0] io_out_bits_payload_manager_xact_id,
  output  io_out_bits_payload_is_builtin_type,
  output [3:0] io_out_bits_payload_g_type,
  output [63:0] io_out_bits_payload_data,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire [1:0] GEN_1;
  wire [1:0] GEN_12;
  wire [1:0] GEN_13;
  wire [1:0] GEN_14;
  wire [1:0] GEN_2;
  wire [1:0] GEN_15;
  wire [1:0] GEN_16;
  wire [1:0] GEN_17;
  wire [2:0] GEN_3;
  wire [2:0] GEN_18;
  wire [2:0] GEN_19;
  wire [2:0] GEN_20;
  wire  GEN_4;
  wire  GEN_21;
  wire  GEN_22;
  wire  GEN_23;
  wire [1:0] GEN_5;
  wire [1:0] GEN_24;
  wire [1:0] GEN_25;
  wire [1:0] GEN_26;
  wire  GEN_6;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_29;
  wire [3:0] GEN_7;
  wire [3:0] GEN_30;
  wire [3:0] GEN_31;
  wire [3:0] GEN_32;
  wire [63:0] GEN_8;
  wire [63:0] GEN_33;
  wire [63:0] GEN_34;
  wire [63:0] GEN_35;
  reg [2:0] T_1100;
  reg [31:0] GEN_47;
  reg [1:0] T_1102;
  reg [31:0] GEN_48;
  wire  T_1104;
  wire [2:0] T_1112_0;
  wire [3:0] GEN_46;
  wire  T_1114;
  wire  T_1115;
  wire  T_1116;
  wire  T_1118;
  wire  T_1119;
  wire [3:0] T_1123;
  wire [2:0] T_1124;
  wire [1:0] GEN_36;
  wire [2:0] GEN_37;
  wire [1:0] GEN_38;
  reg [1:0] lastGrant;
  reg [31:0] GEN_49;
  wire [1:0] GEN_39;
  wire  T_1129;
  wire  T_1131;
  wire  T_1133;
  wire  T_1135;
  wire  T_1136;
  wire  T_1137;
  wire  T_1140;
  wire  T_1141;
  wire  T_1142;
  wire  T_1143;
  wire  T_1144;
  wire  T_1148;
  wire  T_1150;
  wire  T_1152;
  wire  T_1154;
  wire  T_1156;
  wire  T_1158;
  wire  T_1162;
  wire  T_1163;
  wire  T_1164;
  wire  T_1165;
  wire  T_1166;
  wire  T_1168;
  wire  T_1169;
  wire  T_1170;
  wire  T_1172;
  wire  T_1173;
  wire  T_1174;
  wire  T_1176;
  wire  T_1177;
  wire  T_1178;
  wire  T_1180;
  wire  T_1181;
  wire  T_1182;
  wire [1:0] GEN_40;
  wire [1:0] GEN_41;
  wire [1:0] GEN_42;
  wire [1:0] GEN_43;
  wire [1:0] GEN_44;
  wire [1:0] GEN_45;
  assign io_in_0_ready = T_1170;
  assign io_in_1_ready = T_1174;
  assign io_in_2_ready = T_1178;
  assign io_in_3_ready = T_1182;
  assign io_out_valid = GEN_0;
  assign io_out_bits_header_src = GEN_1;
  assign io_out_bits_header_dst = GEN_2;
  assign io_out_bits_payload_addr_beat = GEN_3;
  assign io_out_bits_payload_client_xact_id = GEN_4;
  assign io_out_bits_payload_manager_xact_id = GEN_5;
  assign io_out_bits_payload_is_builtin_type = GEN_6;
  assign io_out_bits_payload_g_type = GEN_7;
  assign io_out_bits_payload_data = GEN_8;
  assign io_chosen = GEN_38;
  assign choice = GEN_45;
  assign GEN_0 = GEN_11;
  assign GEN_9 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_10 = 2'h2 == io_chosen ? io_in_2_valid : GEN_9;
  assign GEN_11 = 2'h3 == io_chosen ? io_in_3_valid : GEN_10;
  assign GEN_1 = GEN_14;
  assign GEN_12 = 2'h1 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_13 = 2'h2 == io_chosen ? io_in_2_bits_header_src : GEN_12;
  assign GEN_14 = 2'h3 == io_chosen ? io_in_3_bits_header_src : GEN_13;
  assign GEN_2 = GEN_17;
  assign GEN_15 = 2'h1 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_16 = 2'h2 == io_chosen ? io_in_2_bits_header_dst : GEN_15;
  assign GEN_17 = 2'h3 == io_chosen ? io_in_3_bits_header_dst : GEN_16;
  assign GEN_3 = GEN_20;
  assign GEN_18 = 2'h1 == io_chosen ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign GEN_19 = 2'h2 == io_chosen ? io_in_2_bits_payload_addr_beat : GEN_18;
  assign GEN_20 = 2'h3 == io_chosen ? io_in_3_bits_payload_addr_beat : GEN_19;
  assign GEN_4 = GEN_23;
  assign GEN_21 = 2'h1 == io_chosen ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign GEN_22 = 2'h2 == io_chosen ? io_in_2_bits_payload_client_xact_id : GEN_21;
  assign GEN_23 = 2'h3 == io_chosen ? io_in_3_bits_payload_client_xact_id : GEN_22;
  assign GEN_5 = GEN_26;
  assign GEN_24 = 2'h1 == io_chosen ? io_in_1_bits_payload_manager_xact_id : io_in_0_bits_payload_manager_xact_id;
  assign GEN_25 = 2'h2 == io_chosen ? io_in_2_bits_payload_manager_xact_id : GEN_24;
  assign GEN_26 = 2'h3 == io_chosen ? io_in_3_bits_payload_manager_xact_id : GEN_25;
  assign GEN_6 = GEN_29;
  assign GEN_27 = 2'h1 == io_chosen ? io_in_1_bits_payload_is_builtin_type : io_in_0_bits_payload_is_builtin_type;
  assign GEN_28 = 2'h2 == io_chosen ? io_in_2_bits_payload_is_builtin_type : GEN_27;
  assign GEN_29 = 2'h3 == io_chosen ? io_in_3_bits_payload_is_builtin_type : GEN_28;
  assign GEN_7 = GEN_32;
  assign GEN_30 = 2'h1 == io_chosen ? io_in_1_bits_payload_g_type : io_in_0_bits_payload_g_type;
  assign GEN_31 = 2'h2 == io_chosen ? io_in_2_bits_payload_g_type : GEN_30;
  assign GEN_32 = 2'h3 == io_chosen ? io_in_3_bits_payload_g_type : GEN_31;
  assign GEN_8 = GEN_35;
  assign GEN_33 = 2'h1 == io_chosen ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign GEN_34 = 2'h2 == io_chosen ? io_in_2_bits_payload_data : GEN_33;
  assign GEN_35 = 2'h3 == io_chosen ? io_in_3_bits_payload_data : GEN_34;
  assign T_1104 = T_1100 != 3'h0;
  assign T_1112_0 = 3'h5;
  assign GEN_46 = {{1'd0}, T_1112_0};
  assign T_1114 = io_out_bits_payload_g_type == GEN_46;
  assign T_1115 = io_out_bits_payload_g_type == 4'h0;
  assign T_1116 = io_out_bits_payload_is_builtin_type ? T_1114 : T_1115;
  assign T_1118 = io_out_ready & io_out_valid;
  assign T_1119 = T_1118 & T_1116;
  assign T_1123 = T_1100 + 3'h1;
  assign T_1124 = T_1123[2:0];
  assign GEN_36 = T_1119 ? io_chosen : T_1102;
  assign GEN_37 = T_1119 ? T_1124 : T_1100;
  assign GEN_38 = T_1104 ? T_1102 : choice;
  assign GEN_39 = T_1118 ? io_chosen : lastGrant;
  assign T_1129 = 2'h1 > lastGrant;
  assign T_1131 = 2'h2 > lastGrant;
  assign T_1133 = 2'h3 > lastGrant;
  assign T_1135 = io_in_1_valid & T_1129;
  assign T_1136 = io_in_2_valid & T_1131;
  assign T_1137 = io_in_3_valid & T_1133;
  assign T_1140 = T_1135 | T_1136;
  assign T_1141 = T_1140 | T_1137;
  assign T_1142 = T_1141 | io_in_0_valid;
  assign T_1143 = T_1142 | io_in_1_valid;
  assign T_1144 = T_1143 | io_in_2_valid;
  assign T_1148 = T_1135 == 1'h0;
  assign T_1150 = T_1140 == 1'h0;
  assign T_1152 = T_1141 == 1'h0;
  assign T_1154 = T_1142 == 1'h0;
  assign T_1156 = T_1143 == 1'h0;
  assign T_1158 = T_1144 == 1'h0;
  assign T_1162 = T_1129 | T_1154;
  assign T_1163 = T_1148 & T_1131;
  assign T_1164 = T_1163 | T_1156;
  assign T_1165 = T_1150 & T_1133;
  assign T_1166 = T_1165 | T_1158;
  assign T_1168 = T_1102 == 2'h0;
  assign T_1169 = T_1104 ? T_1168 : T_1152;
  assign T_1170 = T_1169 & io_out_ready;
  assign T_1172 = T_1102 == 2'h1;
  assign T_1173 = T_1104 ? T_1172 : T_1162;
  assign T_1174 = T_1173 & io_out_ready;
  assign T_1176 = T_1102 == 2'h2;
  assign T_1177 = T_1104 ? T_1176 : T_1164;
  assign T_1178 = T_1177 & io_out_ready;
  assign T_1180 = T_1102 == 2'h3;
  assign T_1181 = T_1104 ? T_1180 : T_1166;
  assign T_1182 = T_1181 & io_out_ready;
  assign GEN_40 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_41 = io_in_1_valid ? 2'h1 : GEN_40;
  assign GEN_42 = io_in_0_valid ? 2'h0 : GEN_41;
  assign GEN_43 = T_1137 ? 2'h3 : GEN_42;
  assign GEN_44 = T_1136 ? 2'h2 : GEN_43;
  assign GEN_45 = T_1135 ? 2'h1 : GEN_44;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_47 = {1{$random}};
  T_1100 = GEN_47[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_48 = {1{$random}};
  T_1102 = GEN_48[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_49 = {1{$random}};
  lastGrant = GEN_49[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1100 <= 3'h0;
    end else begin
      if(T_1119) begin
        T_1100 <= T_1124;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1119) begin
        T_1102 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1118) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module BasicBus_3(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input   io_in_0_bits_payload_client_xact_id,
  input  [1:0] io_in_0_bits_payload_manager_xact_id,
  input   io_in_0_bits_payload_is_builtin_type,
  input  [3:0] io_in_0_bits_payload_g_type,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input   io_in_1_bits_payload_client_xact_id,
  input  [1:0] io_in_1_bits_payload_manager_xact_id,
  input   io_in_1_bits_payload_is_builtin_type,
  input  [3:0] io_in_1_bits_payload_g_type,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input   io_in_2_bits_payload_client_xact_id,
  input  [1:0] io_in_2_bits_payload_manager_xact_id,
  input   io_in_2_bits_payload_is_builtin_type,
  input  [3:0] io_in_2_bits_payload_g_type,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input   io_in_3_bits_payload_client_xact_id,
  input  [1:0] io_in_3_bits_payload_manager_xact_id,
  input   io_in_3_bits_payload_is_builtin_type,
  input  [3:0] io_in_3_bits_payload_g_type,
  input  [63:0] io_in_3_bits_payload_data,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [1:0] io_out_0_bits_header_src,
  output [1:0] io_out_0_bits_header_dst,
  output [2:0] io_out_0_bits_payload_addr_beat,
  output  io_out_0_bits_payload_client_xact_id,
  output [1:0] io_out_0_bits_payload_manager_xact_id,
  output  io_out_0_bits_payload_is_builtin_type,
  output [3:0] io_out_0_bits_payload_g_type,
  output [63:0] io_out_0_bits_payload_data,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [1:0] io_out_1_bits_header_src,
  output [1:0] io_out_1_bits_header_dst,
  output [2:0] io_out_1_bits_payload_addr_beat,
  output  io_out_1_bits_payload_client_xact_id,
  output [1:0] io_out_1_bits_payload_manager_xact_id,
  output  io_out_1_bits_payload_is_builtin_type,
  output [3:0] io_out_1_bits_payload_g_type,
  output [63:0] io_out_1_bits_payload_data,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [1:0] io_out_2_bits_header_src,
  output [1:0] io_out_2_bits_header_dst,
  output [2:0] io_out_2_bits_payload_addr_beat,
  output  io_out_2_bits_payload_client_xact_id,
  output [1:0] io_out_2_bits_payload_manager_xact_id,
  output  io_out_2_bits_payload_is_builtin_type,
  output [3:0] io_out_2_bits_payload_g_type,
  output [63:0] io_out_2_bits_payload_data,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [1:0] io_out_3_bits_header_src,
  output [1:0] io_out_3_bits_header_dst,
  output [2:0] io_out_3_bits_payload_addr_beat,
  output  io_out_3_bits_payload_client_xact_id,
  output [1:0] io_out_3_bits_payload_manager_xact_id,
  output  io_out_3_bits_payload_is_builtin_type,
  output [3:0] io_out_3_bits_payload_g_type,
  output [63:0] io_out_3_bits_payload_data
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_header_src;
  wire [1:0] arb_io_in_0_bits_header_dst;
  wire [2:0] arb_io_in_0_bits_payload_addr_beat;
  wire  arb_io_in_0_bits_payload_client_xact_id;
  wire [1:0] arb_io_in_0_bits_payload_manager_xact_id;
  wire  arb_io_in_0_bits_payload_is_builtin_type;
  wire [3:0] arb_io_in_0_bits_payload_g_type;
  wire [63:0] arb_io_in_0_bits_payload_data;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_header_src;
  wire [1:0] arb_io_in_1_bits_header_dst;
  wire [2:0] arb_io_in_1_bits_payload_addr_beat;
  wire  arb_io_in_1_bits_payload_client_xact_id;
  wire [1:0] arb_io_in_1_bits_payload_manager_xact_id;
  wire  arb_io_in_1_bits_payload_is_builtin_type;
  wire [3:0] arb_io_in_1_bits_payload_g_type;
  wire [63:0] arb_io_in_1_bits_payload_data;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [1:0] arb_io_in_2_bits_header_src;
  wire [1:0] arb_io_in_2_bits_header_dst;
  wire [2:0] arb_io_in_2_bits_payload_addr_beat;
  wire  arb_io_in_2_bits_payload_client_xact_id;
  wire [1:0] arb_io_in_2_bits_payload_manager_xact_id;
  wire  arb_io_in_2_bits_payload_is_builtin_type;
  wire [3:0] arb_io_in_2_bits_payload_g_type;
  wire [63:0] arb_io_in_2_bits_payload_data;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [1:0] arb_io_in_3_bits_header_src;
  wire [1:0] arb_io_in_3_bits_header_dst;
  wire [2:0] arb_io_in_3_bits_payload_addr_beat;
  wire  arb_io_in_3_bits_payload_client_xact_id;
  wire [1:0] arb_io_in_3_bits_payload_manager_xact_id;
  wire  arb_io_in_3_bits_payload_is_builtin_type;
  wire [3:0] arb_io_in_3_bits_payload_g_type;
  wire [63:0] arb_io_in_3_bits_payload_data;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_header_src;
  wire [1:0] arb_io_out_bits_header_dst;
  wire [2:0] arb_io_out_bits_payload_addr_beat;
  wire  arb_io_out_bits_payload_client_xact_id;
  wire [1:0] arb_io_out_bits_payload_manager_xact_id;
  wire  arb_io_out_bits_payload_is_builtin_type;
  wire [3:0] arb_io_out_bits_payload_g_type;
  wire [63:0] arb_io_out_bits_payload_data;
  wire [1:0] arb_io_chosen;
  wire  GEN_0;
  wire  GEN_1;
  wire  GEN_2;
  wire  GEN_3;
  wire  T_1483;
  wire  T_1484;
  wire  T_1486;
  wire  T_1487;
  wire  T_1489;
  wire  T_1490;
  wire  T_1492;
  wire  T_1493;
  LockingRRArbiter_3 arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_beat(arb_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_client_xact_id(arb_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_manager_xact_id(arb_io_in_0_bits_payload_manager_xact_id),
    .io_in_0_bits_payload_is_builtin_type(arb_io_in_0_bits_payload_is_builtin_type),
    .io_in_0_bits_payload_g_type(arb_io_in_0_bits_payload_g_type),
    .io_in_0_bits_payload_data(arb_io_in_0_bits_payload_data),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_beat(arb_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_client_xact_id(arb_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_manager_xact_id(arb_io_in_1_bits_payload_manager_xact_id),
    .io_in_1_bits_payload_is_builtin_type(arb_io_in_1_bits_payload_is_builtin_type),
    .io_in_1_bits_payload_g_type(arb_io_in_1_bits_payload_g_type),
    .io_in_1_bits_payload_data(arb_io_in_1_bits_payload_data),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_beat(arb_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_client_xact_id(arb_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_manager_xact_id(arb_io_in_2_bits_payload_manager_xact_id),
    .io_in_2_bits_payload_is_builtin_type(arb_io_in_2_bits_payload_is_builtin_type),
    .io_in_2_bits_payload_g_type(arb_io_in_2_bits_payload_g_type),
    .io_in_2_bits_payload_data(arb_io_in_2_bits_payload_data),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_beat(arb_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_client_xact_id(arb_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_manager_xact_id(arb_io_in_3_bits_payload_manager_xact_id),
    .io_in_3_bits_payload_is_builtin_type(arb_io_in_3_bits_payload_is_builtin_type),
    .io_in_3_bits_payload_g_type(arb_io_in_3_bits_payload_g_type),
    .io_in_3_bits_payload_data(arb_io_in_3_bits_payload_data),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_addr_beat(arb_io_out_bits_payload_addr_beat),
    .io_out_bits_payload_client_xact_id(arb_io_out_bits_payload_client_xact_id),
    .io_out_bits_payload_manager_xact_id(arb_io_out_bits_payload_manager_xact_id),
    .io_out_bits_payload_is_builtin_type(arb_io_out_bits_payload_is_builtin_type),
    .io_out_bits_payload_g_type(arb_io_out_bits_payload_g_type),
    .io_out_bits_payload_data(arb_io_out_bits_payload_data),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_out_0_valid = T_1484;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_0_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_0_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_0_bits_payload_g_type = arb_io_out_bits_payload_g_type;
  assign io_out_0_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_1_valid = T_1487;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_1_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_1_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_1_bits_payload_g_type = arb_io_out_bits_payload_g_type;
  assign io_out_1_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_2_valid = T_1490;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_2_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_2_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_2_bits_payload_g_type = arb_io_out_bits_payload_g_type;
  assign io_out_2_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_3_valid = T_1493;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_3_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_3_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_3_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_3_bits_payload_g_type = arb_io_out_bits_payload_g_type;
  assign io_out_3_bits_payload_data = arb_io_out_bits_payload_data;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_addr_beat = io_in_0_bits_payload_addr_beat;
  assign arb_io_in_0_bits_payload_client_xact_id = io_in_0_bits_payload_client_xact_id;
  assign arb_io_in_0_bits_payload_manager_xact_id = io_in_0_bits_payload_manager_xact_id;
  assign arb_io_in_0_bits_payload_is_builtin_type = io_in_0_bits_payload_is_builtin_type;
  assign arb_io_in_0_bits_payload_g_type = io_in_0_bits_payload_g_type;
  assign arb_io_in_0_bits_payload_data = io_in_0_bits_payload_data;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_addr_beat = io_in_1_bits_payload_addr_beat;
  assign arb_io_in_1_bits_payload_client_xact_id = io_in_1_bits_payload_client_xact_id;
  assign arb_io_in_1_bits_payload_manager_xact_id = io_in_1_bits_payload_manager_xact_id;
  assign arb_io_in_1_bits_payload_is_builtin_type = io_in_1_bits_payload_is_builtin_type;
  assign arb_io_in_1_bits_payload_g_type = io_in_1_bits_payload_g_type;
  assign arb_io_in_1_bits_payload_data = io_in_1_bits_payload_data;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_addr_beat = io_in_2_bits_payload_addr_beat;
  assign arb_io_in_2_bits_payload_client_xact_id = io_in_2_bits_payload_client_xact_id;
  assign arb_io_in_2_bits_payload_manager_xact_id = io_in_2_bits_payload_manager_xact_id;
  assign arb_io_in_2_bits_payload_is_builtin_type = io_in_2_bits_payload_is_builtin_type;
  assign arb_io_in_2_bits_payload_g_type = io_in_2_bits_payload_g_type;
  assign arb_io_in_2_bits_payload_data = io_in_2_bits_payload_data;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_addr_beat = io_in_3_bits_payload_addr_beat;
  assign arb_io_in_3_bits_payload_client_xact_id = io_in_3_bits_payload_client_xact_id;
  assign arb_io_in_3_bits_payload_manager_xact_id = io_in_3_bits_payload_manager_xact_id;
  assign arb_io_in_3_bits_payload_is_builtin_type = io_in_3_bits_payload_is_builtin_type;
  assign arb_io_in_3_bits_payload_g_type = io_in_3_bits_payload_g_type;
  assign arb_io_in_3_bits_payload_data = io_in_3_bits_payload_data;
  assign arb_io_out_ready = GEN_0;
  assign GEN_0 = GEN_3;
  assign GEN_1 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_2 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_3 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_2;
  assign T_1483 = arb_io_out_bits_header_dst == 2'h0;
  assign T_1484 = arb_io_out_valid & T_1483;
  assign T_1486 = arb_io_out_bits_header_dst == 2'h1;
  assign T_1487 = arb_io_out_valid & T_1486;
  assign T_1489 = arb_io_out_bits_header_dst == 2'h2;
  assign T_1490 = arb_io_out_valid & T_1489;
  assign T_1492 = arb_io_out_bits_header_dst == 2'h3;
  assign T_1493 = arb_io_out_valid & T_1492;
endmodule
module LockingRRArbiter_4(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [1:0] io_in_0_bits_payload_manager_xact_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [1:0] io_in_1_bits_payload_manager_xact_id,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [1:0] io_in_2_bits_payload_manager_xact_id,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [1:0] io_in_3_bits_payload_manager_xact_id,
  input   io_out_ready,
  output  io_out_valid,
  output [1:0] io_out_bits_header_src,
  output [1:0] io_out_bits_header_dst,
  output [1:0] io_out_bits_payload_manager_xact_id,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire [1:0] GEN_1;
  wire [1:0] GEN_7;
  wire [1:0] GEN_8;
  wire [1:0] GEN_9;
  wire [1:0] GEN_2;
  wire [1:0] GEN_10;
  wire [1:0] GEN_11;
  wire [1:0] GEN_12;
  wire [1:0] GEN_3;
  wire [1:0] GEN_13;
  wire [1:0] GEN_14;
  wire [1:0] GEN_15;
  wire  T_930;
  reg [1:0] lastGrant;
  reg [31:0] GEN_23;
  wire [1:0] GEN_16;
  wire  T_933;
  wire  T_935;
  wire  T_937;
  wire  T_939;
  wire  T_940;
  wire  T_941;
  wire  T_944;
  wire  T_945;
  wire  T_946;
  wire  T_947;
  wire  T_948;
  wire  T_952;
  wire  T_954;
  wire  T_956;
  wire  T_958;
  wire  T_960;
  wire  T_962;
  wire  T_966;
  wire  T_967;
  wire  T_968;
  wire  T_969;
  wire  T_970;
  wire  T_971;
  wire  T_972;
  wire  T_973;
  wire  T_974;
  wire [1:0] GEN_17;
  wire [1:0] GEN_18;
  wire [1:0] GEN_19;
  wire [1:0] GEN_20;
  wire [1:0] GEN_21;
  wire [1:0] GEN_22;
  assign io_in_0_ready = T_971;
  assign io_in_1_ready = T_972;
  assign io_in_2_ready = T_973;
  assign io_in_3_ready = T_974;
  assign io_out_valid = GEN_0;
  assign io_out_bits_header_src = GEN_1;
  assign io_out_bits_header_dst = GEN_2;
  assign io_out_bits_payload_manager_xact_id = GEN_3;
  assign io_chosen = choice;
  assign choice = GEN_22;
  assign GEN_0 = GEN_6;
  assign GEN_4 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_5 = 2'h2 == io_chosen ? io_in_2_valid : GEN_4;
  assign GEN_6 = 2'h3 == io_chosen ? io_in_3_valid : GEN_5;
  assign GEN_1 = GEN_9;
  assign GEN_7 = 2'h1 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_8 = 2'h2 == io_chosen ? io_in_2_bits_header_src : GEN_7;
  assign GEN_9 = 2'h3 == io_chosen ? io_in_3_bits_header_src : GEN_8;
  assign GEN_2 = GEN_12;
  assign GEN_10 = 2'h1 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_11 = 2'h2 == io_chosen ? io_in_2_bits_header_dst : GEN_10;
  assign GEN_12 = 2'h3 == io_chosen ? io_in_3_bits_header_dst : GEN_11;
  assign GEN_3 = GEN_15;
  assign GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_payload_manager_xact_id : io_in_0_bits_payload_manager_xact_id;
  assign GEN_14 = 2'h2 == io_chosen ? io_in_2_bits_payload_manager_xact_id : GEN_13;
  assign GEN_15 = 2'h3 == io_chosen ? io_in_3_bits_payload_manager_xact_id : GEN_14;
  assign T_930 = io_out_ready & io_out_valid;
  assign GEN_16 = T_930 ? io_chosen : lastGrant;
  assign T_933 = 2'h1 > lastGrant;
  assign T_935 = 2'h2 > lastGrant;
  assign T_937 = 2'h3 > lastGrant;
  assign T_939 = io_in_1_valid & T_933;
  assign T_940 = io_in_2_valid & T_935;
  assign T_941 = io_in_3_valid & T_937;
  assign T_944 = T_939 | T_940;
  assign T_945 = T_944 | T_941;
  assign T_946 = T_945 | io_in_0_valid;
  assign T_947 = T_946 | io_in_1_valid;
  assign T_948 = T_947 | io_in_2_valid;
  assign T_952 = T_939 == 1'h0;
  assign T_954 = T_944 == 1'h0;
  assign T_956 = T_945 == 1'h0;
  assign T_958 = T_946 == 1'h0;
  assign T_960 = T_947 == 1'h0;
  assign T_962 = T_948 == 1'h0;
  assign T_966 = T_933 | T_958;
  assign T_967 = T_952 & T_935;
  assign T_968 = T_967 | T_960;
  assign T_969 = T_954 & T_937;
  assign T_970 = T_969 | T_962;
  assign T_971 = T_956 & io_out_ready;
  assign T_972 = T_966 & io_out_ready;
  assign T_973 = T_968 & io_out_ready;
  assign T_974 = T_970 & io_out_ready;
  assign GEN_17 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_18 = io_in_1_valid ? 2'h1 : GEN_17;
  assign GEN_19 = io_in_0_valid ? 2'h0 : GEN_18;
  assign GEN_20 = T_941 ? 2'h3 : GEN_19;
  assign GEN_21 = T_940 ? 2'h2 : GEN_20;
  assign GEN_22 = T_939 ? 2'h1 : GEN_21;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_23 = {1{$random}};
  lastGrant = GEN_23[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_930) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module BasicBus_4(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [1:0] io_in_0_bits_header_src,
  input  [1:0] io_in_0_bits_header_dst,
  input  [1:0] io_in_0_bits_payload_manager_xact_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [1:0] io_in_1_bits_header_src,
  input  [1:0] io_in_1_bits_header_dst,
  input  [1:0] io_in_1_bits_payload_manager_xact_id,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [1:0] io_in_2_bits_header_src,
  input  [1:0] io_in_2_bits_header_dst,
  input  [1:0] io_in_2_bits_payload_manager_xact_id,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [1:0] io_in_3_bits_header_src,
  input  [1:0] io_in_3_bits_header_dst,
  input  [1:0] io_in_3_bits_payload_manager_xact_id,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [1:0] io_out_0_bits_header_src,
  output [1:0] io_out_0_bits_header_dst,
  output [1:0] io_out_0_bits_payload_manager_xact_id,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [1:0] io_out_1_bits_header_src,
  output [1:0] io_out_1_bits_header_dst,
  output [1:0] io_out_1_bits_payload_manager_xact_id,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [1:0] io_out_2_bits_header_src,
  output [1:0] io_out_2_bits_header_dst,
  output [1:0] io_out_2_bits_payload_manager_xact_id,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [1:0] io_out_3_bits_header_src,
  output [1:0] io_out_3_bits_header_dst,
  output [1:0] io_out_3_bits_payload_manager_xact_id
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_header_src;
  wire [1:0] arb_io_in_0_bits_header_dst;
  wire [1:0] arb_io_in_0_bits_payload_manager_xact_id;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_header_src;
  wire [1:0] arb_io_in_1_bits_header_dst;
  wire [1:0] arb_io_in_1_bits_payload_manager_xact_id;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [1:0] arb_io_in_2_bits_header_src;
  wire [1:0] arb_io_in_2_bits_header_dst;
  wire [1:0] arb_io_in_2_bits_payload_manager_xact_id;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [1:0] arb_io_in_3_bits_header_src;
  wire [1:0] arb_io_in_3_bits_header_dst;
  wire [1:0] arb_io_in_3_bits_payload_manager_xact_id;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_header_src;
  wire [1:0] arb_io_out_bits_header_dst;
  wire [1:0] arb_io_out_bits_payload_manager_xact_id;
  wire [1:0] arb_io_chosen;
  wire  GEN_0;
  wire  GEN_1;
  wire  GEN_2;
  wire  GEN_3;
  wire  T_1253;
  wire  T_1254;
  wire  T_1256;
  wire  T_1257;
  wire  T_1259;
  wire  T_1260;
  wire  T_1262;
  wire  T_1263;
  LockingRRArbiter_4 arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_manager_xact_id(arb_io_in_0_bits_payload_manager_xact_id),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_manager_xact_id(arb_io_in_1_bits_payload_manager_xact_id),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_manager_xact_id(arb_io_in_2_bits_payload_manager_xact_id),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_manager_xact_id(arb_io_in_3_bits_payload_manager_xact_id),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_manager_xact_id(arb_io_out_bits_payload_manager_xact_id),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_out_0_valid = T_1254;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_1_valid = T_1257;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_2_valid = T_1260;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_3_valid = T_1263;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_manager_xact_id = io_in_0_bits_payload_manager_xact_id;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_manager_xact_id = io_in_1_bits_payload_manager_xact_id;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_manager_xact_id = io_in_2_bits_payload_manager_xact_id;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_manager_xact_id = io_in_3_bits_payload_manager_xact_id;
  assign arb_io_out_ready = GEN_0;
  assign GEN_0 = GEN_3;
  assign GEN_1 = 2'h1 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_2 = 2'h2 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_3 = 2'h3 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_2;
  assign T_1253 = arb_io_out_bits_header_dst == 2'h0;
  assign T_1254 = arb_io_out_valid & T_1253;
  assign T_1256 = arb_io_out_bits_header_dst == 2'h1;
  assign T_1257 = arb_io_out_valid & T_1256;
  assign T_1259 = arb_io_out_bits_header_dst == 2'h2;
  assign T_1260 = arb_io_out_valid & T_1259;
  assign T_1262 = arb_io_out_bits_header_dst == 2'h3;
  assign T_1263 = arb_io_out_valid & T_1262;
endmodule
module PortedTileLinkCrossbar(
  input   clk,
  input   reset,
  output  io_clients_cached_0_acquire_ready,
  input   io_clients_cached_0_acquire_valid,
  input  [25:0] io_clients_cached_0_acquire_bits_addr_block,
  input   io_clients_cached_0_acquire_bits_client_xact_id,
  input  [2:0] io_clients_cached_0_acquire_bits_addr_beat,
  input   io_clients_cached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_clients_cached_0_acquire_bits_a_type,
  input  [11:0] io_clients_cached_0_acquire_bits_union,
  input  [63:0] io_clients_cached_0_acquire_bits_data,
  input   io_clients_cached_0_probe_ready,
  output  io_clients_cached_0_probe_valid,
  output [25:0] io_clients_cached_0_probe_bits_addr_block,
  output [1:0] io_clients_cached_0_probe_bits_p_type,
  output  io_clients_cached_0_release_ready,
  input   io_clients_cached_0_release_valid,
  input  [2:0] io_clients_cached_0_release_bits_addr_beat,
  input  [25:0] io_clients_cached_0_release_bits_addr_block,
  input   io_clients_cached_0_release_bits_client_xact_id,
  input   io_clients_cached_0_release_bits_voluntary,
  input  [2:0] io_clients_cached_0_release_bits_r_type,
  input  [63:0] io_clients_cached_0_release_bits_data,
  input   io_clients_cached_0_grant_ready,
  output  io_clients_cached_0_grant_valid,
  output [2:0] io_clients_cached_0_grant_bits_addr_beat,
  output  io_clients_cached_0_grant_bits_client_xact_id,
  output [1:0] io_clients_cached_0_grant_bits_manager_xact_id,
  output  io_clients_cached_0_grant_bits_is_builtin_type,
  output [3:0] io_clients_cached_0_grant_bits_g_type,
  output [63:0] io_clients_cached_0_grant_bits_data,
  output  io_clients_cached_0_grant_bits_manager_id,
  output  io_clients_cached_0_finish_ready,
  input   io_clients_cached_0_finish_valid,
  input  [1:0] io_clients_cached_0_finish_bits_manager_xact_id,
  input   io_clients_cached_0_finish_bits_manager_id,
  output  io_clients_uncached_0_acquire_ready,
  input   io_clients_uncached_0_acquire_valid,
  input  [25:0] io_clients_uncached_0_acquire_bits_addr_block,
  input   io_clients_uncached_0_acquire_bits_client_xact_id,
  input  [2:0] io_clients_uncached_0_acquire_bits_addr_beat,
  input   io_clients_uncached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_clients_uncached_0_acquire_bits_a_type,
  input  [11:0] io_clients_uncached_0_acquire_bits_union,
  input  [63:0] io_clients_uncached_0_acquire_bits_data,
  input   io_clients_uncached_0_grant_ready,
  output  io_clients_uncached_0_grant_valid,
  output [2:0] io_clients_uncached_0_grant_bits_addr_beat,
  output  io_clients_uncached_0_grant_bits_client_xact_id,
  output [1:0] io_clients_uncached_0_grant_bits_manager_xact_id,
  output  io_clients_uncached_0_grant_bits_is_builtin_type,
  output [3:0] io_clients_uncached_0_grant_bits_g_type,
  output [63:0] io_clients_uncached_0_grant_bits_data,
  input   io_managers_0_acquire_ready,
  output  io_managers_0_acquire_valid,
  output [25:0] io_managers_0_acquire_bits_addr_block,
  output  io_managers_0_acquire_bits_client_xact_id,
  output [2:0] io_managers_0_acquire_bits_addr_beat,
  output  io_managers_0_acquire_bits_is_builtin_type,
  output [2:0] io_managers_0_acquire_bits_a_type,
  output [11:0] io_managers_0_acquire_bits_union,
  output [63:0] io_managers_0_acquire_bits_data,
  output  io_managers_0_acquire_bits_client_id,
  output  io_managers_0_grant_ready,
  input   io_managers_0_grant_valid,
  input  [2:0] io_managers_0_grant_bits_addr_beat,
  input   io_managers_0_grant_bits_client_xact_id,
  input  [1:0] io_managers_0_grant_bits_manager_xact_id,
  input   io_managers_0_grant_bits_is_builtin_type,
  input  [3:0] io_managers_0_grant_bits_g_type,
  input  [63:0] io_managers_0_grant_bits_data,
  input   io_managers_0_grant_bits_client_id,
  input   io_managers_0_finish_ready,
  output  io_managers_0_finish_valid,
  output [1:0] io_managers_0_finish_bits_manager_xact_id,
  output  io_managers_0_probe_ready,
  input   io_managers_0_probe_valid,
  input  [25:0] io_managers_0_probe_bits_addr_block,
  input  [1:0] io_managers_0_probe_bits_p_type,
  input   io_managers_0_probe_bits_client_id,
  input   io_managers_0_release_ready,
  output  io_managers_0_release_valid,
  output [2:0] io_managers_0_release_bits_addr_beat,
  output [25:0] io_managers_0_release_bits_addr_block,
  output  io_managers_0_release_bits_client_xact_id,
  output  io_managers_0_release_bits_voluntary,
  output [2:0] io_managers_0_release_bits_r_type,
  output [63:0] io_managers_0_release_bits_data,
  output  io_managers_0_release_bits_client_id,
  input   io_managers_1_acquire_ready,
  output  io_managers_1_acquire_valid,
  output [25:0] io_managers_1_acquire_bits_addr_block,
  output  io_managers_1_acquire_bits_client_xact_id,
  output [2:0] io_managers_1_acquire_bits_addr_beat,
  output  io_managers_1_acquire_bits_is_builtin_type,
  output [2:0] io_managers_1_acquire_bits_a_type,
  output [11:0] io_managers_1_acquire_bits_union,
  output [63:0] io_managers_1_acquire_bits_data,
  output  io_managers_1_acquire_bits_client_id,
  output  io_managers_1_grant_ready,
  input   io_managers_1_grant_valid,
  input  [2:0] io_managers_1_grant_bits_addr_beat,
  input   io_managers_1_grant_bits_client_xact_id,
  input  [1:0] io_managers_1_grant_bits_manager_xact_id,
  input   io_managers_1_grant_bits_is_builtin_type,
  input  [3:0] io_managers_1_grant_bits_g_type,
  input  [63:0] io_managers_1_grant_bits_data,
  input   io_managers_1_grant_bits_client_id,
  input   io_managers_1_finish_ready,
  output  io_managers_1_finish_valid,
  output [1:0] io_managers_1_finish_bits_manager_xact_id,
  output  io_managers_1_probe_ready,
  input   io_managers_1_probe_valid,
  input  [25:0] io_managers_1_probe_bits_addr_block,
  input  [1:0] io_managers_1_probe_bits_p_type,
  input   io_managers_1_probe_bits_client_id,
  input   io_managers_1_release_ready,
  output  io_managers_1_release_valid,
  output [2:0] io_managers_1_release_bits_addr_beat,
  output [25:0] io_managers_1_release_bits_addr_block,
  output  io_managers_1_release_bits_client_xact_id,
  output  io_managers_1_release_bits_voluntary,
  output [2:0] io_managers_1_release_bits_r_type,
  output [63:0] io_managers_1_release_bits_data,
  output  io_managers_1_release_bits_client_id
);
  wire  TileLinkEnqueuer_4_clk;
  wire  TileLinkEnqueuer_4_reset;
  wire  TileLinkEnqueuer_4_io_client_acquire_ready;
  wire  TileLinkEnqueuer_4_io_client_acquire_valid;
  wire [1:0] TileLinkEnqueuer_4_io_client_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_client_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_block;
  wire  TileLinkEnqueuer_4_io_client_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_4_io_client_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_4_io_client_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_4_io_client_grant_ready;
  wire  TileLinkEnqueuer_4_io_client_grant_valid;
  wire [1:0] TileLinkEnqueuer_4_io_client_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_client_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_4_io_client_grant_bits_payload_client_xact_id;
  wire [1:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_4_io_client_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_4_io_client_grant_bits_payload_data;
  wire  TileLinkEnqueuer_4_io_client_finish_ready;
  wire  TileLinkEnqueuer_4_io_client_finish_valid;
  wire [1:0] TileLinkEnqueuer_4_io_client_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_client_finish_bits_header_dst;
  wire [1:0] TileLinkEnqueuer_4_io_client_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_4_io_client_probe_ready;
  wire  TileLinkEnqueuer_4_io_client_probe_valid;
  wire [1:0] TileLinkEnqueuer_4_io_client_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_client_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_4_io_client_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_io_client_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_4_io_client_release_ready;
  wire  TileLinkEnqueuer_4_io_client_release_valid;
  wire [1:0] TileLinkEnqueuer_4_io_client_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_client_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_io_client_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_4_io_client_release_bits_payload_addr_block;
  wire  TileLinkEnqueuer_4_io_client_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_4_io_client_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_4_io_client_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_4_io_client_release_bits_payload_data;
  wire  TileLinkEnqueuer_4_io_manager_acquire_ready;
  wire  TileLinkEnqueuer_4_io_manager_acquire_valid;
  wire [1:0] TileLinkEnqueuer_4_io_manager_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_manager_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_block;
  wire  TileLinkEnqueuer_4_io_manager_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_4_io_manager_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_4_io_manager_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_4_io_manager_grant_ready;
  wire  TileLinkEnqueuer_4_io_manager_grant_valid;
  wire [1:0] TileLinkEnqueuer_4_io_manager_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_manager_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_io_manager_grant_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_4_io_manager_grant_bits_payload_client_xact_id;
  wire [1:0] TileLinkEnqueuer_4_io_manager_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_4_io_manager_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_4_io_manager_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_4_io_manager_grant_bits_payload_data;
  wire  TileLinkEnqueuer_4_io_manager_finish_ready;
  wire  TileLinkEnqueuer_4_io_manager_finish_valid;
  wire [1:0] TileLinkEnqueuer_4_io_manager_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_manager_finish_bits_header_dst;
  wire [1:0] TileLinkEnqueuer_4_io_manager_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_4_io_manager_probe_ready;
  wire  TileLinkEnqueuer_4_io_manager_probe_valid;
  wire [1:0] TileLinkEnqueuer_4_io_manager_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_manager_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_4_io_manager_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_io_manager_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_4_io_manager_release_ready;
  wire  TileLinkEnqueuer_4_io_manager_release_valid;
  wire [1:0] TileLinkEnqueuer_4_io_manager_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_4_io_manager_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_block;
  wire  TileLinkEnqueuer_4_io_manager_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_4_io_manager_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_4_io_manager_release_bits_payload_data;
  wire  ClientTileLinkNetworkPort_1_clk;
  wire  ClientTileLinkNetworkPort_1_reset;
  wire  ClientTileLinkNetworkPort_1_io_client_acquire_ready;
  wire  ClientTileLinkNetworkPort_1_io_client_acquire_valid;
  wire [25:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_block;
  wire  ClientTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat;
  wire  ClientTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_a_type;
  wire [11:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_union;
  wire [63:0] ClientTileLinkNetworkPort_1_io_client_acquire_bits_data;
  wire  ClientTileLinkNetworkPort_1_io_client_probe_ready;
  wire  ClientTileLinkNetworkPort_1_io_client_probe_valid;
  wire [25:0] ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type;
  wire  ClientTileLinkNetworkPort_1_io_client_release_ready;
  wire  ClientTileLinkNetworkPort_1_io_client_release_valid;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_release_bits_addr_beat;
  wire [25:0] ClientTileLinkNetworkPort_1_io_client_release_bits_addr_block;
  wire  ClientTileLinkNetworkPort_1_io_client_release_bits_client_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_client_release_bits_voluntary;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_release_bits_r_type;
  wire [63:0] ClientTileLinkNetworkPort_1_io_client_release_bits_data;
  wire  ClientTileLinkNetworkPort_1_io_client_grant_ready;
  wire  ClientTileLinkNetworkPort_1_io_client_grant_valid;
  wire [2:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  wire  ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  wire [1:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  wire [63:0] ClientTileLinkNetworkPort_1_io_client_grant_bits_data;
  wire  ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_id;
  wire  ClientTileLinkNetworkPort_1_io_client_finish_ready;
  wire  ClientTileLinkNetworkPort_1_io_client_finish_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_id;
  wire  ClientTileLinkNetworkPort_1_io_network_acquire_ready;
  wire  ClientTileLinkNetworkPort_1_io_network_acquire_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst;
  wire [25:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block;
  wire  ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat;
  wire  ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type;
  wire [11:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union;
  wire [63:0] ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data;
  wire  ClientTileLinkNetworkPort_1_io_network_grant_ready;
  wire  ClientTileLinkNetworkPort_1_io_network_grant_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_header_src;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_header_dst;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat;
  wire  ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type;
  wire [3:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type;
  wire [63:0] ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_data;
  wire  ClientTileLinkNetworkPort_1_io_network_finish_ready;
  wire  ClientTileLinkNetworkPort_1_io_network_finish_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_network_probe_ready;
  wire  ClientTileLinkNetworkPort_1_io_network_probe_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_probe_bits_header_src;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_probe_bits_header_dst;
  wire [25:0] ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type;
  wire  ClientTileLinkNetworkPort_1_io_network_release_ready;
  wire  ClientTileLinkNetworkPort_1_io_network_release_valid;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_header_src;
  wire [1:0] ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat;
  wire [25:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block;
  wire  ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id;
  wire  ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary;
  wire [2:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type;
  wire [63:0] ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_clk;
  wire  TileLinkEnqueuer_1_1_reset;
  wire  TileLinkEnqueuer_1_1_io_client_acquire_ready;
  wire  TileLinkEnqueuer_1_1_io_client_acquire_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_block;
  wire  TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_io_client_grant_ready;
  wire  TileLinkEnqueuer_1_1_io_client_grant_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_grant_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_1_1_io_client_grant_bits_payload_client_xact_id;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_1_1_io_client_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_1_1_io_client_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_1_1_io_client_grant_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_io_client_finish_ready;
  wire  TileLinkEnqueuer_1_1_io_client_finish_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_finish_bits_header_dst;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_1_1_io_client_probe_ready;
  wire  TileLinkEnqueuer_1_1_io_client_probe_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_1_1_io_client_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_1_1_io_client_release_ready;
  wire  TileLinkEnqueuer_1_1_io_client_release_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_client_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_block;
  wire  TileLinkEnqueuer_1_1_io_client_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_1_1_io_client_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_1_1_io_client_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_1_1_io_client_release_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_io_manager_acquire_ready;
  wire  TileLinkEnqueuer_1_1_io_manager_acquire_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_block;
  wire  TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_io_manager_grant_ready;
  wire  TileLinkEnqueuer_1_1_io_manager_grant_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_client_xact_id;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_data;
  wire  TileLinkEnqueuer_1_1_io_manager_finish_ready;
  wire  TileLinkEnqueuer_1_1_io_manager_finish_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_finish_bits_header_dst;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_1_1_io_manager_probe_ready;
  wire  TileLinkEnqueuer_1_1_io_manager_probe_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_1_1_io_manager_release_ready;
  wire  TileLinkEnqueuer_1_1_io_manager_release_valid;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_1_1_io_manager_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_block;
  wire  TileLinkEnqueuer_1_1_io_manager_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_1_1_io_manager_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_1_1_io_manager_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_1_1_io_manager_release_bits_payload_data;
  wire  ClientUncachedTileLinkNetworkPort_1_clk;
  wire  ClientUncachedTileLinkNetworkPort_1_reset;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_acquire_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_acquire_valid;
  wire [25:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_block;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_data;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_grant_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_grant_valid;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_data;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_acquire_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_acquire_valid;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_src;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_dst;
  wire [25:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type;
  wire [11:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_union;
  wire [63:0] ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_data;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_grant_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_grant_valid;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_src;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_dst;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type;
  wire [63:0] ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_data;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_finish_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_finish_valid;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_src;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_dst;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_probe_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_probe_valid;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_src;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_dst;
  wire [25:0] ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_release_ready;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_release_valid;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_src;
  wire [1:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_dst;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat;
  wire [25:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary;
  wire [2:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_r_type;
  wire [63:0] ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_2_clk;
  wire  ManagerTileLinkNetworkPort_2_reset;
  wire  ManagerTileLinkNetworkPort_2_io_manager_acquire_ready;
  wire  ManagerTileLinkNetworkPort_2_io_manager_acquire_valid;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_block;
  wire  ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_beat;
  wire  ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_is_builtin_type;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_a_type;
  wire [11:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_union;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_data;
  wire  ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_grant_ready;
  wire  ManagerTileLinkNetworkPort_2_io_manager_grant_valid;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_grant_bits_addr_beat;
  wire  ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_xact_id;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_manager_grant_bits_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_grant_bits_is_builtin_type;
  wire [3:0] ManagerTileLinkNetworkPort_2_io_manager_grant_bits_g_type;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_manager_grant_bits_data;
  wire  ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_finish_ready;
  wire  ManagerTileLinkNetworkPort_2_io_manager_finish_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_manager_finish_bits_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_probe_ready;
  wire  ManagerTileLinkNetworkPort_2_io_manager_probe_valid;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_manager_probe_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_manager_probe_bits_p_type;
  wire  ManagerTileLinkNetworkPort_2_io_manager_probe_bits_client_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_release_ready;
  wire  ManagerTileLinkNetworkPort_2_io_manager_release_valid;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_beat;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_block;
  wire  ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_manager_release_bits_voluntary;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_manager_release_bits_r_type;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_manager_release_bits_data;
  wire  ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_id;
  wire  ManagerTileLinkNetworkPort_2_io_network_acquire_ready;
  wire  ManagerTileLinkNetworkPort_2_io_network_acquire_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_dst;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block;
  wire  ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat;
  wire  ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type;
  wire [11:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_union;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_2_io_network_grant_ready;
  wire  ManagerTileLinkNetworkPort_2_io_network_grant_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_addr_beat;
  wire  ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_client_xact_id;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_is_builtin_type;
  wire [3:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_g_type;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_2_io_network_finish_ready;
  wire  ManagerTileLinkNetworkPort_2_io_network_finish_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_dst;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_network_probe_ready;
  wire  ManagerTileLinkNetworkPort_2_io_network_probe_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_dst;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_p_type;
  wire  ManagerTileLinkNetworkPort_2_io_network_release_ready;
  wire  ManagerTileLinkNetworkPort_2_io_network_release_valid;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat;
  wire [25:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block;
  wire  ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id;
  wire  ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary;
  wire [2:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_r_type;
  wire [63:0] ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_clk;
  wire  TileLinkEnqueuer_2_1_reset;
  wire  TileLinkEnqueuer_2_1_io_client_acquire_ready;
  wire  TileLinkEnqueuer_2_1_io_client_acquire_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_block;
  wire  TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_io_client_grant_ready;
  wire  TileLinkEnqueuer_2_1_io_client_grant_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_grant_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_2_1_io_client_grant_bits_payload_client_xact_id;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_2_1_io_client_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_2_1_io_client_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_2_1_io_client_grant_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_io_client_finish_ready;
  wire  TileLinkEnqueuer_2_1_io_client_finish_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_finish_bits_header_dst;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_2_1_io_client_probe_ready;
  wire  TileLinkEnqueuer_2_1_io_client_probe_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_2_1_io_client_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_2_1_io_client_release_ready;
  wire  TileLinkEnqueuer_2_1_io_client_release_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_client_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_block;
  wire  TileLinkEnqueuer_2_1_io_client_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_2_1_io_client_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_2_1_io_client_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_2_1_io_client_release_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_io_manager_acquire_ready;
  wire  TileLinkEnqueuer_2_1_io_manager_acquire_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_block;
  wire  TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_io_manager_grant_ready;
  wire  TileLinkEnqueuer_2_1_io_manager_grant_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_client_xact_id;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_data;
  wire  TileLinkEnqueuer_2_1_io_manager_finish_ready;
  wire  TileLinkEnqueuer_2_1_io_manager_finish_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_finish_bits_header_dst;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_2_1_io_manager_probe_ready;
  wire  TileLinkEnqueuer_2_1_io_manager_probe_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_2_1_io_manager_release_ready;
  wire  TileLinkEnqueuer_2_1_io_manager_release_valid;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_2_1_io_manager_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_block;
  wire  TileLinkEnqueuer_2_1_io_manager_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_2_1_io_manager_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_2_1_io_manager_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_2_1_io_manager_release_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_1_1_clk;
  wire  ManagerTileLinkNetworkPort_1_1_reset;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_acquire_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_acquire_valid;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_block;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_beat;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_is_builtin_type;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_a_type;
  wire [11:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_union;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_data;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_grant_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_grant_valid;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_addr_beat;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_xact_id;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_is_builtin_type;
  wire [3:0] ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_g_type;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_data;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_finish_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_finish_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_manager_finish_bits_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_probe_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_probe_valid;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_p_type;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_client_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_release_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_release_valid;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_beat;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_block;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_voluntary;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_r_type;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_data;
  wire  ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_acquire_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_acquire_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_dst;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_block;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_beat;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_is_builtin_type;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_a_type;
  wire [11:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_union;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_grant_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_grant_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_addr_beat;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_client_xact_id;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_is_builtin_type;
  wire [3:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_g_type;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_finish_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_finish_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_dst;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_payload_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_probe_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_probe_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_dst;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_p_type;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_release_ready;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_release_valid;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_src;
  wire [1:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_beat;
  wire [25:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_block;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_client_xact_id;
  wire  ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_voluntary;
  wire [2:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_r_type;
  wire [63:0] ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_clk;
  wire  TileLinkEnqueuer_3_1_reset;
  wire  TileLinkEnqueuer_3_1_io_client_acquire_ready;
  wire  TileLinkEnqueuer_3_1_io_client_acquire_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_block;
  wire  TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_io_client_grant_ready;
  wire  TileLinkEnqueuer_3_1_io_client_grant_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_grant_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_3_1_io_client_grant_bits_payload_client_xact_id;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_3_1_io_client_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_3_1_io_client_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_3_1_io_client_grant_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_io_client_finish_ready;
  wire  TileLinkEnqueuer_3_1_io_client_finish_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_finish_bits_header_dst;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_3_1_io_client_probe_ready;
  wire  TileLinkEnqueuer_3_1_io_client_probe_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_3_1_io_client_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_3_1_io_client_release_ready;
  wire  TileLinkEnqueuer_3_1_io_client_release_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_client_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_block;
  wire  TileLinkEnqueuer_3_1_io_client_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_3_1_io_client_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_3_1_io_client_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_3_1_io_client_release_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_io_manager_acquire_ready;
  wire  TileLinkEnqueuer_3_1_io_manager_acquire_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_block;
  wire  TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_io_manager_grant_ready;
  wire  TileLinkEnqueuer_3_1_io_manager_grant_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_client_xact_id;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_data;
  wire  TileLinkEnqueuer_3_1_io_manager_finish_ready;
  wire  TileLinkEnqueuer_3_1_io_manager_finish_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_finish_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_finish_bits_header_dst;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_3_1_io_manager_probe_ready;
  wire  TileLinkEnqueuer_3_1_io_manager_probe_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_probe_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_3_1_io_manager_release_ready;
  wire  TileLinkEnqueuer_3_1_io_manager_release_valid;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_release_bits_header_src;
  wire [1:0] TileLinkEnqueuer_3_1_io_manager_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_block;
  wire  TileLinkEnqueuer_3_1_io_manager_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_3_1_io_manager_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_3_1_io_manager_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_3_1_io_manager_release_bits_payload_data;
  wire  acqNet_clk;
  wire  acqNet_reset;
  wire  acqNet_io_in_0_ready;
  wire  acqNet_io_in_0_valid;
  wire [1:0] acqNet_io_in_0_bits_header_src;
  wire [1:0] acqNet_io_in_0_bits_header_dst;
  wire [25:0] acqNet_io_in_0_bits_payload_addr_block;
  wire  acqNet_io_in_0_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_in_0_bits_payload_addr_beat;
  wire  acqNet_io_in_0_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_in_0_bits_payload_a_type;
  wire [11:0] acqNet_io_in_0_bits_payload_union;
  wire [63:0] acqNet_io_in_0_bits_payload_data;
  wire  acqNet_io_in_1_ready;
  wire  acqNet_io_in_1_valid;
  wire [1:0] acqNet_io_in_1_bits_header_src;
  wire [1:0] acqNet_io_in_1_bits_header_dst;
  wire [25:0] acqNet_io_in_1_bits_payload_addr_block;
  wire  acqNet_io_in_1_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_in_1_bits_payload_addr_beat;
  wire  acqNet_io_in_1_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_in_1_bits_payload_a_type;
  wire [11:0] acqNet_io_in_1_bits_payload_union;
  wire [63:0] acqNet_io_in_1_bits_payload_data;
  wire  acqNet_io_in_2_ready;
  wire  acqNet_io_in_2_valid;
  wire [1:0] acqNet_io_in_2_bits_header_src;
  wire [1:0] acqNet_io_in_2_bits_header_dst;
  wire [25:0] acqNet_io_in_2_bits_payload_addr_block;
  wire  acqNet_io_in_2_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_in_2_bits_payload_addr_beat;
  wire  acqNet_io_in_2_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_in_2_bits_payload_a_type;
  wire [11:0] acqNet_io_in_2_bits_payload_union;
  wire [63:0] acqNet_io_in_2_bits_payload_data;
  wire  acqNet_io_in_3_ready;
  wire  acqNet_io_in_3_valid;
  wire [1:0] acqNet_io_in_3_bits_header_src;
  wire [1:0] acqNet_io_in_3_bits_header_dst;
  wire [25:0] acqNet_io_in_3_bits_payload_addr_block;
  wire  acqNet_io_in_3_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_in_3_bits_payload_addr_beat;
  wire  acqNet_io_in_3_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_in_3_bits_payload_a_type;
  wire [11:0] acqNet_io_in_3_bits_payload_union;
  wire [63:0] acqNet_io_in_3_bits_payload_data;
  wire  acqNet_io_out_0_ready;
  wire  acqNet_io_out_0_valid;
  wire [1:0] acqNet_io_out_0_bits_header_src;
  wire [1:0] acqNet_io_out_0_bits_header_dst;
  wire [25:0] acqNet_io_out_0_bits_payload_addr_block;
  wire  acqNet_io_out_0_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_out_0_bits_payload_addr_beat;
  wire  acqNet_io_out_0_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_out_0_bits_payload_a_type;
  wire [11:0] acqNet_io_out_0_bits_payload_union;
  wire [63:0] acqNet_io_out_0_bits_payload_data;
  wire  acqNet_io_out_1_ready;
  wire  acqNet_io_out_1_valid;
  wire [1:0] acqNet_io_out_1_bits_header_src;
  wire [1:0] acqNet_io_out_1_bits_header_dst;
  wire [25:0] acqNet_io_out_1_bits_payload_addr_block;
  wire  acqNet_io_out_1_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_out_1_bits_payload_addr_beat;
  wire  acqNet_io_out_1_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_out_1_bits_payload_a_type;
  wire [11:0] acqNet_io_out_1_bits_payload_union;
  wire [63:0] acqNet_io_out_1_bits_payload_data;
  wire  acqNet_io_out_2_ready;
  wire  acqNet_io_out_2_valid;
  wire [1:0] acqNet_io_out_2_bits_header_src;
  wire [1:0] acqNet_io_out_2_bits_header_dst;
  wire [25:0] acqNet_io_out_2_bits_payload_addr_block;
  wire  acqNet_io_out_2_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_out_2_bits_payload_addr_beat;
  wire  acqNet_io_out_2_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_out_2_bits_payload_a_type;
  wire [11:0] acqNet_io_out_2_bits_payload_union;
  wire [63:0] acqNet_io_out_2_bits_payload_data;
  wire  acqNet_io_out_3_ready;
  wire  acqNet_io_out_3_valid;
  wire [1:0] acqNet_io_out_3_bits_header_src;
  wire [1:0] acqNet_io_out_3_bits_header_dst;
  wire [25:0] acqNet_io_out_3_bits_payload_addr_block;
  wire  acqNet_io_out_3_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_out_3_bits_payload_addr_beat;
  wire  acqNet_io_out_3_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_out_3_bits_payload_a_type;
  wire [11:0] acqNet_io_out_3_bits_payload_union;
  wire [63:0] acqNet_io_out_3_bits_payload_data;
  wire  relNet_clk;
  wire  relNet_reset;
  wire  relNet_io_in_0_ready;
  wire  relNet_io_in_0_valid;
  wire [1:0] relNet_io_in_0_bits_header_src;
  wire [1:0] relNet_io_in_0_bits_header_dst;
  wire [2:0] relNet_io_in_0_bits_payload_addr_beat;
  wire [25:0] relNet_io_in_0_bits_payload_addr_block;
  wire  relNet_io_in_0_bits_payload_client_xact_id;
  wire  relNet_io_in_0_bits_payload_voluntary;
  wire [2:0] relNet_io_in_0_bits_payload_r_type;
  wire [63:0] relNet_io_in_0_bits_payload_data;
  wire  relNet_io_in_1_ready;
  wire  relNet_io_in_1_valid;
  wire [1:0] relNet_io_in_1_bits_header_src;
  wire [1:0] relNet_io_in_1_bits_header_dst;
  wire [2:0] relNet_io_in_1_bits_payload_addr_beat;
  wire [25:0] relNet_io_in_1_bits_payload_addr_block;
  wire  relNet_io_in_1_bits_payload_client_xact_id;
  wire  relNet_io_in_1_bits_payload_voluntary;
  wire [2:0] relNet_io_in_1_bits_payload_r_type;
  wire [63:0] relNet_io_in_1_bits_payload_data;
  wire  relNet_io_in_2_ready;
  wire  relNet_io_in_2_valid;
  wire [1:0] relNet_io_in_2_bits_header_src;
  wire [1:0] relNet_io_in_2_bits_header_dst;
  wire [2:0] relNet_io_in_2_bits_payload_addr_beat;
  wire [25:0] relNet_io_in_2_bits_payload_addr_block;
  wire  relNet_io_in_2_bits_payload_client_xact_id;
  wire  relNet_io_in_2_bits_payload_voluntary;
  wire [2:0] relNet_io_in_2_bits_payload_r_type;
  wire [63:0] relNet_io_in_2_bits_payload_data;
  wire  relNet_io_in_3_ready;
  wire  relNet_io_in_3_valid;
  wire [1:0] relNet_io_in_3_bits_header_src;
  wire [1:0] relNet_io_in_3_bits_header_dst;
  wire [2:0] relNet_io_in_3_bits_payload_addr_beat;
  wire [25:0] relNet_io_in_3_bits_payload_addr_block;
  wire  relNet_io_in_3_bits_payload_client_xact_id;
  wire  relNet_io_in_3_bits_payload_voluntary;
  wire [2:0] relNet_io_in_3_bits_payload_r_type;
  wire [63:0] relNet_io_in_3_bits_payload_data;
  wire  relNet_io_out_0_ready;
  wire  relNet_io_out_0_valid;
  wire [1:0] relNet_io_out_0_bits_header_src;
  wire [1:0] relNet_io_out_0_bits_header_dst;
  wire [2:0] relNet_io_out_0_bits_payload_addr_beat;
  wire [25:0] relNet_io_out_0_bits_payload_addr_block;
  wire  relNet_io_out_0_bits_payload_client_xact_id;
  wire  relNet_io_out_0_bits_payload_voluntary;
  wire [2:0] relNet_io_out_0_bits_payload_r_type;
  wire [63:0] relNet_io_out_0_bits_payload_data;
  wire  relNet_io_out_1_ready;
  wire  relNet_io_out_1_valid;
  wire [1:0] relNet_io_out_1_bits_header_src;
  wire [1:0] relNet_io_out_1_bits_header_dst;
  wire [2:0] relNet_io_out_1_bits_payload_addr_beat;
  wire [25:0] relNet_io_out_1_bits_payload_addr_block;
  wire  relNet_io_out_1_bits_payload_client_xact_id;
  wire  relNet_io_out_1_bits_payload_voluntary;
  wire [2:0] relNet_io_out_1_bits_payload_r_type;
  wire [63:0] relNet_io_out_1_bits_payload_data;
  wire  relNet_io_out_2_ready;
  wire  relNet_io_out_2_valid;
  wire [1:0] relNet_io_out_2_bits_header_src;
  wire [1:0] relNet_io_out_2_bits_header_dst;
  wire [2:0] relNet_io_out_2_bits_payload_addr_beat;
  wire [25:0] relNet_io_out_2_bits_payload_addr_block;
  wire  relNet_io_out_2_bits_payload_client_xact_id;
  wire  relNet_io_out_2_bits_payload_voluntary;
  wire [2:0] relNet_io_out_2_bits_payload_r_type;
  wire [63:0] relNet_io_out_2_bits_payload_data;
  wire  relNet_io_out_3_ready;
  wire  relNet_io_out_3_valid;
  wire [1:0] relNet_io_out_3_bits_header_src;
  wire [1:0] relNet_io_out_3_bits_header_dst;
  wire [2:0] relNet_io_out_3_bits_payload_addr_beat;
  wire [25:0] relNet_io_out_3_bits_payload_addr_block;
  wire  relNet_io_out_3_bits_payload_client_xact_id;
  wire  relNet_io_out_3_bits_payload_voluntary;
  wire [2:0] relNet_io_out_3_bits_payload_r_type;
  wire [63:0] relNet_io_out_3_bits_payload_data;
  wire  prbNet_clk;
  wire  prbNet_reset;
  wire  prbNet_io_in_0_ready;
  wire  prbNet_io_in_0_valid;
  wire [1:0] prbNet_io_in_0_bits_header_src;
  wire [1:0] prbNet_io_in_0_bits_header_dst;
  wire [25:0] prbNet_io_in_0_bits_payload_addr_block;
  wire [1:0] prbNet_io_in_0_bits_payload_p_type;
  wire  prbNet_io_in_1_ready;
  wire  prbNet_io_in_1_valid;
  wire [1:0] prbNet_io_in_1_bits_header_src;
  wire [1:0] prbNet_io_in_1_bits_header_dst;
  wire [25:0] prbNet_io_in_1_bits_payload_addr_block;
  wire [1:0] prbNet_io_in_1_bits_payload_p_type;
  wire  prbNet_io_in_2_ready;
  wire  prbNet_io_in_2_valid;
  wire [1:0] prbNet_io_in_2_bits_header_src;
  wire [1:0] prbNet_io_in_2_bits_header_dst;
  wire [25:0] prbNet_io_in_2_bits_payload_addr_block;
  wire [1:0] prbNet_io_in_2_bits_payload_p_type;
  wire  prbNet_io_in_3_ready;
  wire  prbNet_io_in_3_valid;
  wire [1:0] prbNet_io_in_3_bits_header_src;
  wire [1:0] prbNet_io_in_3_bits_header_dst;
  wire [25:0] prbNet_io_in_3_bits_payload_addr_block;
  wire [1:0] prbNet_io_in_3_bits_payload_p_type;
  wire  prbNet_io_out_0_ready;
  wire  prbNet_io_out_0_valid;
  wire [1:0] prbNet_io_out_0_bits_header_src;
  wire [1:0] prbNet_io_out_0_bits_header_dst;
  wire [25:0] prbNet_io_out_0_bits_payload_addr_block;
  wire [1:0] prbNet_io_out_0_bits_payload_p_type;
  wire  prbNet_io_out_1_ready;
  wire  prbNet_io_out_1_valid;
  wire [1:0] prbNet_io_out_1_bits_header_src;
  wire [1:0] prbNet_io_out_1_bits_header_dst;
  wire [25:0] prbNet_io_out_1_bits_payload_addr_block;
  wire [1:0] prbNet_io_out_1_bits_payload_p_type;
  wire  prbNet_io_out_2_ready;
  wire  prbNet_io_out_2_valid;
  wire [1:0] prbNet_io_out_2_bits_header_src;
  wire [1:0] prbNet_io_out_2_bits_header_dst;
  wire [25:0] prbNet_io_out_2_bits_payload_addr_block;
  wire [1:0] prbNet_io_out_2_bits_payload_p_type;
  wire  prbNet_io_out_3_ready;
  wire  prbNet_io_out_3_valid;
  wire [1:0] prbNet_io_out_3_bits_header_src;
  wire [1:0] prbNet_io_out_3_bits_header_dst;
  wire [25:0] prbNet_io_out_3_bits_payload_addr_block;
  wire [1:0] prbNet_io_out_3_bits_payload_p_type;
  wire  gntNet_clk;
  wire  gntNet_reset;
  wire  gntNet_io_in_0_ready;
  wire  gntNet_io_in_0_valid;
  wire [1:0] gntNet_io_in_0_bits_header_src;
  wire [1:0] gntNet_io_in_0_bits_header_dst;
  wire [2:0] gntNet_io_in_0_bits_payload_addr_beat;
  wire  gntNet_io_in_0_bits_payload_client_xact_id;
  wire [1:0] gntNet_io_in_0_bits_payload_manager_xact_id;
  wire  gntNet_io_in_0_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_in_0_bits_payload_g_type;
  wire [63:0] gntNet_io_in_0_bits_payload_data;
  wire  gntNet_io_in_1_ready;
  wire  gntNet_io_in_1_valid;
  wire [1:0] gntNet_io_in_1_bits_header_src;
  wire [1:0] gntNet_io_in_1_bits_header_dst;
  wire [2:0] gntNet_io_in_1_bits_payload_addr_beat;
  wire  gntNet_io_in_1_bits_payload_client_xact_id;
  wire [1:0] gntNet_io_in_1_bits_payload_manager_xact_id;
  wire  gntNet_io_in_1_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_in_1_bits_payload_g_type;
  wire [63:0] gntNet_io_in_1_bits_payload_data;
  wire  gntNet_io_in_2_ready;
  wire  gntNet_io_in_2_valid;
  wire [1:0] gntNet_io_in_2_bits_header_src;
  wire [1:0] gntNet_io_in_2_bits_header_dst;
  wire [2:0] gntNet_io_in_2_bits_payload_addr_beat;
  wire  gntNet_io_in_2_bits_payload_client_xact_id;
  wire [1:0] gntNet_io_in_2_bits_payload_manager_xact_id;
  wire  gntNet_io_in_2_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_in_2_bits_payload_g_type;
  wire [63:0] gntNet_io_in_2_bits_payload_data;
  wire  gntNet_io_in_3_ready;
  wire  gntNet_io_in_3_valid;
  wire [1:0] gntNet_io_in_3_bits_header_src;
  wire [1:0] gntNet_io_in_3_bits_header_dst;
  wire [2:0] gntNet_io_in_3_bits_payload_addr_beat;
  wire  gntNet_io_in_3_bits_payload_client_xact_id;
  wire [1:0] gntNet_io_in_3_bits_payload_manager_xact_id;
  wire  gntNet_io_in_3_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_in_3_bits_payload_g_type;
  wire [63:0] gntNet_io_in_3_bits_payload_data;
  wire  gntNet_io_out_0_ready;
  wire  gntNet_io_out_0_valid;
  wire [1:0] gntNet_io_out_0_bits_header_src;
  wire [1:0] gntNet_io_out_0_bits_header_dst;
  wire [2:0] gntNet_io_out_0_bits_payload_addr_beat;
  wire  gntNet_io_out_0_bits_payload_client_xact_id;
  wire [1:0] gntNet_io_out_0_bits_payload_manager_xact_id;
  wire  gntNet_io_out_0_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_out_0_bits_payload_g_type;
  wire [63:0] gntNet_io_out_0_bits_payload_data;
  wire  gntNet_io_out_1_ready;
  wire  gntNet_io_out_1_valid;
  wire [1:0] gntNet_io_out_1_bits_header_src;
  wire [1:0] gntNet_io_out_1_bits_header_dst;
  wire [2:0] gntNet_io_out_1_bits_payload_addr_beat;
  wire  gntNet_io_out_1_bits_payload_client_xact_id;
  wire [1:0] gntNet_io_out_1_bits_payload_manager_xact_id;
  wire  gntNet_io_out_1_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_out_1_bits_payload_g_type;
  wire [63:0] gntNet_io_out_1_bits_payload_data;
  wire  gntNet_io_out_2_ready;
  wire  gntNet_io_out_2_valid;
  wire [1:0] gntNet_io_out_2_bits_header_src;
  wire [1:0] gntNet_io_out_2_bits_header_dst;
  wire [2:0] gntNet_io_out_2_bits_payload_addr_beat;
  wire  gntNet_io_out_2_bits_payload_client_xact_id;
  wire [1:0] gntNet_io_out_2_bits_payload_manager_xact_id;
  wire  gntNet_io_out_2_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_out_2_bits_payload_g_type;
  wire [63:0] gntNet_io_out_2_bits_payload_data;
  wire  gntNet_io_out_3_ready;
  wire  gntNet_io_out_3_valid;
  wire [1:0] gntNet_io_out_3_bits_header_src;
  wire [1:0] gntNet_io_out_3_bits_header_dst;
  wire [2:0] gntNet_io_out_3_bits_payload_addr_beat;
  wire  gntNet_io_out_3_bits_payload_client_xact_id;
  wire [1:0] gntNet_io_out_3_bits_payload_manager_xact_id;
  wire  gntNet_io_out_3_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_out_3_bits_payload_g_type;
  wire [63:0] gntNet_io_out_3_bits_payload_data;
  wire  ackNet_clk;
  wire  ackNet_reset;
  wire  ackNet_io_in_0_ready;
  wire  ackNet_io_in_0_valid;
  wire [1:0] ackNet_io_in_0_bits_header_src;
  wire [1:0] ackNet_io_in_0_bits_header_dst;
  wire [1:0] ackNet_io_in_0_bits_payload_manager_xact_id;
  wire  ackNet_io_in_1_ready;
  wire  ackNet_io_in_1_valid;
  wire [1:0] ackNet_io_in_1_bits_header_src;
  wire [1:0] ackNet_io_in_1_bits_header_dst;
  wire [1:0] ackNet_io_in_1_bits_payload_manager_xact_id;
  wire  ackNet_io_in_2_ready;
  wire  ackNet_io_in_2_valid;
  wire [1:0] ackNet_io_in_2_bits_header_src;
  wire [1:0] ackNet_io_in_2_bits_header_dst;
  wire [1:0] ackNet_io_in_2_bits_payload_manager_xact_id;
  wire  ackNet_io_in_3_ready;
  wire  ackNet_io_in_3_valid;
  wire [1:0] ackNet_io_in_3_bits_header_src;
  wire [1:0] ackNet_io_in_3_bits_header_dst;
  wire [1:0] ackNet_io_in_3_bits_payload_manager_xact_id;
  wire  ackNet_io_out_0_ready;
  wire  ackNet_io_out_0_valid;
  wire [1:0] ackNet_io_out_0_bits_header_src;
  wire [1:0] ackNet_io_out_0_bits_header_dst;
  wire [1:0] ackNet_io_out_0_bits_payload_manager_xact_id;
  wire  ackNet_io_out_1_ready;
  wire  ackNet_io_out_1_valid;
  wire [1:0] ackNet_io_out_1_bits_header_src;
  wire [1:0] ackNet_io_out_1_bits_header_dst;
  wire [1:0] ackNet_io_out_1_bits_payload_manager_xact_id;
  wire  ackNet_io_out_2_ready;
  wire  ackNet_io_out_2_valid;
  wire [1:0] ackNet_io_out_2_bits_header_src;
  wire [1:0] ackNet_io_out_2_bits_header_dst;
  wire [1:0] ackNet_io_out_2_bits_payload_manager_xact_id;
  wire  ackNet_io_out_3_ready;
  wire  ackNet_io_out_3_valid;
  wire [1:0] ackNet_io_out_3_bits_header_src;
  wire [1:0] ackNet_io_out_3_bits_header_dst;
  wire [1:0] ackNet_io_out_3_bits_payload_manager_xact_id;
  wire  T_12724_ready;
  wire  T_12724_valid;
  wire [1:0] T_12724_bits_header_src;
  wire [1:0] T_12724_bits_header_dst;
  wire [25:0] T_12724_bits_payload_addr_block;
  wire  T_12724_bits_payload_client_xact_id;
  wire [2:0] T_12724_bits_payload_addr_beat;
  wire  T_12724_bits_payload_is_builtin_type;
  wire [2:0] T_12724_bits_payload_a_type;
  wire [11:0] T_12724_bits_payload_union;
  wire [63:0] T_12724_bits_payload_data;
  wire [2:0] T_12952;
  wire [1:0] T_12953;
  wire  T_13294_ready;
  wire  T_13294_valid;
  wire [1:0] T_13294_bits_header_src;
  wire [1:0] T_13294_bits_header_dst;
  wire [25:0] T_13294_bits_payload_addr_block;
  wire  T_13294_bits_payload_client_xact_id;
  wire [2:0] T_13294_bits_payload_addr_beat;
  wire  T_13294_bits_payload_is_builtin_type;
  wire [2:0] T_13294_bits_payload_a_type;
  wire [11:0] T_13294_bits_payload_union;
  wire [63:0] T_13294_bits_payload_data;
  wire [2:0] T_13522;
  wire [1:0] T_13523;
  wire  T_13624_ready;
  wire  T_13624_valid;
  wire [1:0] T_13624_bits_header_src;
  wire [1:0] T_13624_bits_header_dst;
  wire [25:0] T_13624_bits_payload_addr_block;
  wire  T_13624_bits_payload_client_xact_id;
  wire [2:0] T_13624_bits_payload_addr_beat;
  wire  T_13624_bits_payload_is_builtin_type;
  wire [2:0] T_13624_bits_payload_a_type;
  wire [11:0] T_13624_bits_payload_union;
  wire [63:0] T_13624_bits_payload_data;
  wire [2:0] T_13692;
  wire [1:0] T_13693;
  wire  T_13794_ready;
  wire  T_13794_valid;
  wire [1:0] T_13794_bits_header_src;
  wire [1:0] T_13794_bits_header_dst;
  wire [25:0] T_13794_bits_payload_addr_block;
  wire  T_13794_bits_payload_client_xact_id;
  wire [2:0] T_13794_bits_payload_addr_beat;
  wire  T_13794_bits_payload_is_builtin_type;
  wire [2:0] T_13794_bits_payload_a_type;
  wire [11:0] T_13794_bits_payload_union;
  wire [63:0] T_13794_bits_payload_data;
  wire [2:0] T_13862;
  wire [1:0] T_13863;
  wire  T_14201_ready;
  wire  T_14201_valid;
  wire [1:0] T_14201_bits_header_src;
  wire [1:0] T_14201_bits_header_dst;
  wire [2:0] T_14201_bits_payload_addr_beat;
  wire [25:0] T_14201_bits_payload_addr_block;
  wire  T_14201_bits_payload_client_xact_id;
  wire  T_14201_bits_payload_voluntary;
  wire [2:0] T_14201_bits_payload_r_type;
  wire [63:0] T_14201_bits_payload_data;
  wire [2:0] T_14427;
  wire [1:0] T_14428;
  wire  T_14766_ready;
  wire  T_14766_valid;
  wire [1:0] T_14766_bits_header_src;
  wire [1:0] T_14766_bits_header_dst;
  wire [2:0] T_14766_bits_payload_addr_beat;
  wire [25:0] T_14766_bits_payload_addr_block;
  wire  T_14766_bits_payload_client_xact_id;
  wire  T_14766_bits_payload_voluntary;
  wire [2:0] T_14766_bits_payload_r_type;
  wire [63:0] T_14766_bits_payload_data;
  wire [2:0] T_14992;
  wire [1:0] T_14993;
  wire  T_15091_ready;
  wire  T_15091_valid;
  wire [1:0] T_15091_bits_header_src;
  wire [1:0] T_15091_bits_header_dst;
  wire [2:0] T_15091_bits_payload_addr_beat;
  wire [25:0] T_15091_bits_payload_addr_block;
  wire  T_15091_bits_payload_client_xact_id;
  wire  T_15091_bits_payload_voluntary;
  wire [2:0] T_15091_bits_payload_r_type;
  wire [63:0] T_15091_bits_payload_data;
  wire [2:0] T_15157;
  wire [1:0] T_15158;
  wire  T_15256_ready;
  wire  T_15256_valid;
  wire [1:0] T_15256_bits_header_src;
  wire [1:0] T_15256_bits_header_dst;
  wire [2:0] T_15256_bits_payload_addr_beat;
  wire [25:0] T_15256_bits_payload_addr_block;
  wire  T_15256_bits_payload_client_xact_id;
  wire  T_15256_bits_payload_voluntary;
  wire [2:0] T_15256_bits_payload_r_type;
  wire [63:0] T_15256_bits_payload_data;
  wire [2:0] T_15322;
  wire [1:0] T_15323;
  wire  T_15409_ready;
  wire  T_15409_valid;
  wire [1:0] T_15409_bits_header_src;
  wire [1:0] T_15409_bits_header_dst;
  wire [25:0] T_15409_bits_payload_addr_block;
  wire [1:0] T_15409_bits_payload_p_type;
  wire [2:0] T_15467;
  wire [1:0] T_15468;
  wire  T_15554_ready;
  wire  T_15554_valid;
  wire [1:0] T_15554_bits_header_src;
  wire [1:0] T_15554_bits_header_dst;
  wire [25:0] T_15554_bits_payload_addr_block;
  wire [1:0] T_15554_bits_payload_p_type;
  wire [2:0] T_15612;
  wire [1:0] T_15613;
  wire  T_15939_ready;
  wire  T_15939_valid;
  wire [1:0] T_15939_bits_header_src;
  wire [1:0] T_15939_bits_header_dst;
  wire [25:0] T_15939_bits_payload_addr_block;
  wire [1:0] T_15939_bits_payload_p_type;
  wire [2:0] T_16157;
  wire [1:0] T_16158;
  wire  T_16484_ready;
  wire  T_16484_valid;
  wire [1:0] T_16484_bits_header_src;
  wire [1:0] T_16484_bits_header_dst;
  wire [25:0] T_16484_bits_payload_addr_block;
  wire [1:0] T_16484_bits_payload_p_type;
  wire [2:0] T_16702;
  wire [1:0] T_16703;
  wire  T_16801_ready;
  wire  T_16801_valid;
  wire [1:0] T_16801_bits_header_src;
  wire [1:0] T_16801_bits_header_dst;
  wire [2:0] T_16801_bits_payload_addr_beat;
  wire  T_16801_bits_payload_client_xact_id;
  wire [1:0] T_16801_bits_payload_manager_xact_id;
  wire  T_16801_bits_payload_is_builtin_type;
  wire [3:0] T_16801_bits_payload_g_type;
  wire [63:0] T_16801_bits_payload_data;
  wire [2:0] T_16867;
  wire [1:0] T_16868;
  wire  T_16966_ready;
  wire  T_16966_valid;
  wire [1:0] T_16966_bits_header_src;
  wire [1:0] T_16966_bits_header_dst;
  wire [2:0] T_16966_bits_payload_addr_beat;
  wire  T_16966_bits_payload_client_xact_id;
  wire [1:0] T_16966_bits_payload_manager_xact_id;
  wire  T_16966_bits_payload_is_builtin_type;
  wire [3:0] T_16966_bits_payload_g_type;
  wire [63:0] T_16966_bits_payload_data;
  wire [2:0] T_17032;
  wire [1:0] T_17033;
  wire  T_17371_ready;
  wire  T_17371_valid;
  wire [1:0] T_17371_bits_header_src;
  wire [1:0] T_17371_bits_header_dst;
  wire [2:0] T_17371_bits_payload_addr_beat;
  wire  T_17371_bits_payload_client_xact_id;
  wire [1:0] T_17371_bits_payload_manager_xact_id;
  wire  T_17371_bits_payload_is_builtin_type;
  wire [3:0] T_17371_bits_payload_g_type;
  wire [63:0] T_17371_bits_payload_data;
  wire [2:0] T_17597;
  wire [1:0] T_17598;
  wire  T_17936_ready;
  wire  T_17936_valid;
  wire [1:0] T_17936_bits_header_src;
  wire [1:0] T_17936_bits_header_dst;
  wire [2:0] T_17936_bits_payload_addr_beat;
  wire  T_17936_bits_payload_client_xact_id;
  wire [1:0] T_17936_bits_payload_manager_xact_id;
  wire  T_17936_bits_payload_is_builtin_type;
  wire [3:0] T_17936_bits_payload_g_type;
  wire [63:0] T_17936_bits_payload_data;
  wire [2:0] T_18162;
  wire [1:0] T_18163;
  wire  T_18486_ready;
  wire  T_18486_valid;
  wire [1:0] T_18486_bits_header_src;
  wire [1:0] T_18486_bits_header_dst;
  wire [1:0] T_18486_bits_payload_manager_xact_id;
  wire [2:0] T_18702;
  wire [1:0] T_18703;
  wire  T_19026_ready;
  wire  T_19026_valid;
  wire [1:0] T_19026_bits_header_src;
  wire [1:0] T_19026_bits_header_dst;
  wire [1:0] T_19026_bits_payload_manager_xact_id;
  wire [2:0] T_19242;
  wire [1:0] T_19243;
  wire  T_19326_ready;
  wire  T_19326_valid;
  wire [1:0] T_19326_bits_header_src;
  wire [1:0] T_19326_bits_header_dst;
  wire [1:0] T_19326_bits_payload_manager_xact_id;
  wire [2:0] T_19382;
  wire [1:0] T_19383;
  wire  T_19466_ready;
  wire  T_19466_valid;
  wire [1:0] T_19466_bits_header_src;
  wire [1:0] T_19466_bits_header_dst;
  wire [1:0] T_19466_bits_payload_manager_xact_id;
  wire [2:0] T_19522;
  wire [1:0] T_19523;
  reg [1:0] GEN_0;
  reg [31:0] GEN_64;
  reg [1:0] GEN_1;
  reg [31:0] GEN_65;
  reg [25:0] GEN_2;
  reg [31:0] GEN_66;
  reg  GEN_3;
  reg [31:0] GEN_67;
  reg [2:0] GEN_4;
  reg [31:0] GEN_68;
  reg  GEN_5;
  reg [31:0] GEN_69;
  reg [2:0] GEN_6;
  reg [31:0] GEN_70;
  reg [11:0] GEN_7;
  reg [31:0] GEN_71;
  reg [63:0] GEN_8;
  reg [63:0] GEN_72;
  reg [1:0] GEN_9;
  reg [31:0] GEN_73;
  reg [1:0] GEN_10;
  reg [31:0] GEN_74;
  reg [25:0] GEN_11;
  reg [31:0] GEN_75;
  reg  GEN_12;
  reg [31:0] GEN_76;
  reg [2:0] GEN_13;
  reg [31:0] GEN_77;
  reg  GEN_14;
  reg [31:0] GEN_78;
  reg [2:0] GEN_15;
  reg [31:0] GEN_79;
  reg [11:0] GEN_16;
  reg [31:0] GEN_80;
  reg [63:0] GEN_17;
  reg [63:0] GEN_81;
  reg [1:0] GEN_18;
  reg [31:0] GEN_82;
  reg [1:0] GEN_19;
  reg [31:0] GEN_83;
  reg [2:0] GEN_20;
  reg [31:0] GEN_84;
  reg [25:0] GEN_21;
  reg [31:0] GEN_85;
  reg  GEN_22;
  reg [31:0] GEN_86;
  reg  GEN_23;
  reg [31:0] GEN_87;
  reg [2:0] GEN_24;
  reg [31:0] GEN_88;
  reg [63:0] GEN_25;
  reg [63:0] GEN_89;
  reg [1:0] GEN_26;
  reg [31:0] GEN_90;
  reg [1:0] GEN_27;
  reg [31:0] GEN_91;
  reg [2:0] GEN_28;
  reg [31:0] GEN_92;
  reg [25:0] GEN_29;
  reg [31:0] GEN_93;
  reg  GEN_30;
  reg [31:0] GEN_94;
  reg  GEN_31;
  reg [31:0] GEN_95;
  reg [2:0] GEN_32;
  reg [31:0] GEN_96;
  reg [63:0] GEN_33;
  reg [63:0] GEN_97;
  reg [1:0] GEN_34;
  reg [31:0] GEN_98;
  reg [1:0] GEN_35;
  reg [31:0] GEN_99;
  reg [25:0] GEN_36;
  reg [31:0] GEN_100;
  reg [1:0] GEN_37;
  reg [31:0] GEN_101;
  reg [1:0] GEN_38;
  reg [31:0] GEN_102;
  reg [1:0] GEN_39;
  reg [31:0] GEN_103;
  reg [25:0] GEN_40;
  reg [31:0] GEN_104;
  reg [1:0] GEN_41;
  reg [31:0] GEN_105;
  reg [1:0] GEN_42;
  reg [31:0] GEN_106;
  reg [1:0] GEN_43;
  reg [31:0] GEN_107;
  reg [2:0] GEN_44;
  reg [31:0] GEN_108;
  reg  GEN_45;
  reg [31:0] GEN_109;
  reg [1:0] GEN_46;
  reg [31:0] GEN_110;
  reg  GEN_47;
  reg [31:0] GEN_111;
  reg [3:0] GEN_48;
  reg [31:0] GEN_112;
  reg [63:0] GEN_49;
  reg [63:0] GEN_113;
  reg [1:0] GEN_50;
  reg [31:0] GEN_114;
  reg [1:0] GEN_51;
  reg [31:0] GEN_115;
  reg [2:0] GEN_52;
  reg [31:0] GEN_116;
  reg  GEN_53;
  reg [31:0] GEN_117;
  reg [1:0] GEN_54;
  reg [31:0] GEN_118;
  reg  GEN_55;
  reg [31:0] GEN_119;
  reg [3:0] GEN_56;
  reg [31:0] GEN_120;
  reg [63:0] GEN_57;
  reg [63:0] GEN_121;
  reg [1:0] GEN_58;
  reg [31:0] GEN_122;
  reg [1:0] GEN_59;
  reg [31:0] GEN_123;
  reg [1:0] GEN_60;
  reg [31:0] GEN_124;
  reg [1:0] GEN_61;
  reg [31:0] GEN_125;
  reg [1:0] GEN_62;
  reg [31:0] GEN_126;
  reg [1:0] GEN_63;
  reg [31:0] GEN_127;
  TileLinkEnqueuer TileLinkEnqueuer_4 (
    .clk(TileLinkEnqueuer_4_clk),
    .reset(TileLinkEnqueuer_4_reset),
    .io_client_acquire_ready(TileLinkEnqueuer_4_io_client_acquire_ready),
    .io_client_acquire_valid(TileLinkEnqueuer_4_io_client_acquire_valid),
    .io_client_acquire_bits_header_src(TileLinkEnqueuer_4_io_client_acquire_bits_header_src),
    .io_client_acquire_bits_header_dst(TileLinkEnqueuer_4_io_client_acquire_bits_header_dst),
    .io_client_acquire_bits_payload_addr_block(TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_block),
    .io_client_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_client_acquire_bits_payload_client_xact_id),
    .io_client_acquire_bits_payload_addr_beat(TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_beat),
    .io_client_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_4_io_client_acquire_bits_payload_is_builtin_type),
    .io_client_acquire_bits_payload_a_type(TileLinkEnqueuer_4_io_client_acquire_bits_payload_a_type),
    .io_client_acquire_bits_payload_union(TileLinkEnqueuer_4_io_client_acquire_bits_payload_union),
    .io_client_acquire_bits_payload_data(TileLinkEnqueuer_4_io_client_acquire_bits_payload_data),
    .io_client_grant_ready(TileLinkEnqueuer_4_io_client_grant_ready),
    .io_client_grant_valid(TileLinkEnqueuer_4_io_client_grant_valid),
    .io_client_grant_bits_header_src(TileLinkEnqueuer_4_io_client_grant_bits_header_src),
    .io_client_grant_bits_header_dst(TileLinkEnqueuer_4_io_client_grant_bits_header_dst),
    .io_client_grant_bits_payload_addr_beat(TileLinkEnqueuer_4_io_client_grant_bits_payload_addr_beat),
    .io_client_grant_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_client_grant_bits_payload_client_xact_id),
    .io_client_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_4_io_client_grant_bits_payload_manager_xact_id),
    .io_client_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_4_io_client_grant_bits_payload_is_builtin_type),
    .io_client_grant_bits_payload_g_type(TileLinkEnqueuer_4_io_client_grant_bits_payload_g_type),
    .io_client_grant_bits_payload_data(TileLinkEnqueuer_4_io_client_grant_bits_payload_data),
    .io_client_finish_ready(TileLinkEnqueuer_4_io_client_finish_ready),
    .io_client_finish_valid(TileLinkEnqueuer_4_io_client_finish_valid),
    .io_client_finish_bits_header_src(TileLinkEnqueuer_4_io_client_finish_bits_header_src),
    .io_client_finish_bits_header_dst(TileLinkEnqueuer_4_io_client_finish_bits_header_dst),
    .io_client_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_4_io_client_finish_bits_payload_manager_xact_id),
    .io_client_probe_ready(TileLinkEnqueuer_4_io_client_probe_ready),
    .io_client_probe_valid(TileLinkEnqueuer_4_io_client_probe_valid),
    .io_client_probe_bits_header_src(TileLinkEnqueuer_4_io_client_probe_bits_header_src),
    .io_client_probe_bits_header_dst(TileLinkEnqueuer_4_io_client_probe_bits_header_dst),
    .io_client_probe_bits_payload_addr_block(TileLinkEnqueuer_4_io_client_probe_bits_payload_addr_block),
    .io_client_probe_bits_payload_p_type(TileLinkEnqueuer_4_io_client_probe_bits_payload_p_type),
    .io_client_release_ready(TileLinkEnqueuer_4_io_client_release_ready),
    .io_client_release_valid(TileLinkEnqueuer_4_io_client_release_valid),
    .io_client_release_bits_header_src(TileLinkEnqueuer_4_io_client_release_bits_header_src),
    .io_client_release_bits_header_dst(TileLinkEnqueuer_4_io_client_release_bits_header_dst),
    .io_client_release_bits_payload_addr_beat(TileLinkEnqueuer_4_io_client_release_bits_payload_addr_beat),
    .io_client_release_bits_payload_addr_block(TileLinkEnqueuer_4_io_client_release_bits_payload_addr_block),
    .io_client_release_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_client_release_bits_payload_client_xact_id),
    .io_client_release_bits_payload_voluntary(TileLinkEnqueuer_4_io_client_release_bits_payload_voluntary),
    .io_client_release_bits_payload_r_type(TileLinkEnqueuer_4_io_client_release_bits_payload_r_type),
    .io_client_release_bits_payload_data(TileLinkEnqueuer_4_io_client_release_bits_payload_data),
    .io_manager_acquire_ready(TileLinkEnqueuer_4_io_manager_acquire_ready),
    .io_manager_acquire_valid(TileLinkEnqueuer_4_io_manager_acquire_valid),
    .io_manager_acquire_bits_header_src(TileLinkEnqueuer_4_io_manager_acquire_bits_header_src),
    .io_manager_acquire_bits_header_dst(TileLinkEnqueuer_4_io_manager_acquire_bits_header_dst),
    .io_manager_acquire_bits_payload_addr_block(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_block),
    .io_manager_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_client_xact_id),
    .io_manager_acquire_bits_payload_addr_beat(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_beat),
    .io_manager_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_is_builtin_type),
    .io_manager_acquire_bits_payload_a_type(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_a_type),
    .io_manager_acquire_bits_payload_union(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_union),
    .io_manager_acquire_bits_payload_data(TileLinkEnqueuer_4_io_manager_acquire_bits_payload_data),
    .io_manager_grant_ready(TileLinkEnqueuer_4_io_manager_grant_ready),
    .io_manager_grant_valid(TileLinkEnqueuer_4_io_manager_grant_valid),
    .io_manager_grant_bits_header_src(TileLinkEnqueuer_4_io_manager_grant_bits_header_src),
    .io_manager_grant_bits_header_dst(TileLinkEnqueuer_4_io_manager_grant_bits_header_dst),
    .io_manager_grant_bits_payload_addr_beat(TileLinkEnqueuer_4_io_manager_grant_bits_payload_addr_beat),
    .io_manager_grant_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_manager_grant_bits_payload_client_xact_id),
    .io_manager_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_4_io_manager_grant_bits_payload_manager_xact_id),
    .io_manager_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_4_io_manager_grant_bits_payload_is_builtin_type),
    .io_manager_grant_bits_payload_g_type(TileLinkEnqueuer_4_io_manager_grant_bits_payload_g_type),
    .io_manager_grant_bits_payload_data(TileLinkEnqueuer_4_io_manager_grant_bits_payload_data),
    .io_manager_finish_ready(TileLinkEnqueuer_4_io_manager_finish_ready),
    .io_manager_finish_valid(TileLinkEnqueuer_4_io_manager_finish_valid),
    .io_manager_finish_bits_header_src(TileLinkEnqueuer_4_io_manager_finish_bits_header_src),
    .io_manager_finish_bits_header_dst(TileLinkEnqueuer_4_io_manager_finish_bits_header_dst),
    .io_manager_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_4_io_manager_finish_bits_payload_manager_xact_id),
    .io_manager_probe_ready(TileLinkEnqueuer_4_io_manager_probe_ready),
    .io_manager_probe_valid(TileLinkEnqueuer_4_io_manager_probe_valid),
    .io_manager_probe_bits_header_src(TileLinkEnqueuer_4_io_manager_probe_bits_header_src),
    .io_manager_probe_bits_header_dst(TileLinkEnqueuer_4_io_manager_probe_bits_header_dst),
    .io_manager_probe_bits_payload_addr_block(TileLinkEnqueuer_4_io_manager_probe_bits_payload_addr_block),
    .io_manager_probe_bits_payload_p_type(TileLinkEnqueuer_4_io_manager_probe_bits_payload_p_type),
    .io_manager_release_ready(TileLinkEnqueuer_4_io_manager_release_ready),
    .io_manager_release_valid(TileLinkEnqueuer_4_io_manager_release_valid),
    .io_manager_release_bits_header_src(TileLinkEnqueuer_4_io_manager_release_bits_header_src),
    .io_manager_release_bits_header_dst(TileLinkEnqueuer_4_io_manager_release_bits_header_dst),
    .io_manager_release_bits_payload_addr_beat(TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_beat),
    .io_manager_release_bits_payload_addr_block(TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_block),
    .io_manager_release_bits_payload_client_xact_id(TileLinkEnqueuer_4_io_manager_release_bits_payload_client_xact_id),
    .io_manager_release_bits_payload_voluntary(TileLinkEnqueuer_4_io_manager_release_bits_payload_voluntary),
    .io_manager_release_bits_payload_r_type(TileLinkEnqueuer_4_io_manager_release_bits_payload_r_type),
    .io_manager_release_bits_payload_data(TileLinkEnqueuer_4_io_manager_release_bits_payload_data)
  );
  ClientTileLinkNetworkPort ClientTileLinkNetworkPort_1 (
    .clk(ClientTileLinkNetworkPort_1_clk),
    .reset(ClientTileLinkNetworkPort_1_reset),
    .io_client_acquire_ready(ClientTileLinkNetworkPort_1_io_client_acquire_ready),
    .io_client_acquire_valid(ClientTileLinkNetworkPort_1_io_client_acquire_valid),
    .io_client_acquire_bits_addr_block(ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_block),
    .io_client_acquire_bits_client_xact_id(ClientTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id),
    .io_client_acquire_bits_addr_beat(ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat),
    .io_client_acquire_bits_is_builtin_type(ClientTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type),
    .io_client_acquire_bits_a_type(ClientTileLinkNetworkPort_1_io_client_acquire_bits_a_type),
    .io_client_acquire_bits_union(ClientTileLinkNetworkPort_1_io_client_acquire_bits_union),
    .io_client_acquire_bits_data(ClientTileLinkNetworkPort_1_io_client_acquire_bits_data),
    .io_client_probe_ready(ClientTileLinkNetworkPort_1_io_client_probe_ready),
    .io_client_probe_valid(ClientTileLinkNetworkPort_1_io_client_probe_valid),
    .io_client_probe_bits_addr_block(ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block),
    .io_client_probe_bits_p_type(ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type),
    .io_client_release_ready(ClientTileLinkNetworkPort_1_io_client_release_ready),
    .io_client_release_valid(ClientTileLinkNetworkPort_1_io_client_release_valid),
    .io_client_release_bits_addr_beat(ClientTileLinkNetworkPort_1_io_client_release_bits_addr_beat),
    .io_client_release_bits_addr_block(ClientTileLinkNetworkPort_1_io_client_release_bits_addr_block),
    .io_client_release_bits_client_xact_id(ClientTileLinkNetworkPort_1_io_client_release_bits_client_xact_id),
    .io_client_release_bits_voluntary(ClientTileLinkNetworkPort_1_io_client_release_bits_voluntary),
    .io_client_release_bits_r_type(ClientTileLinkNetworkPort_1_io_client_release_bits_r_type),
    .io_client_release_bits_data(ClientTileLinkNetworkPort_1_io_client_release_bits_data),
    .io_client_grant_ready(ClientTileLinkNetworkPort_1_io_client_grant_ready),
    .io_client_grant_valid(ClientTileLinkNetworkPort_1_io_client_grant_valid),
    .io_client_grant_bits_addr_beat(ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat),
    .io_client_grant_bits_client_xact_id(ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id),
    .io_client_grant_bits_manager_xact_id(ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id),
    .io_client_grant_bits_is_builtin_type(ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type),
    .io_client_grant_bits_g_type(ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type),
    .io_client_grant_bits_data(ClientTileLinkNetworkPort_1_io_client_grant_bits_data),
    .io_client_grant_bits_manager_id(ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_id),
    .io_client_finish_ready(ClientTileLinkNetworkPort_1_io_client_finish_ready),
    .io_client_finish_valid(ClientTileLinkNetworkPort_1_io_client_finish_valid),
    .io_client_finish_bits_manager_xact_id(ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_xact_id),
    .io_client_finish_bits_manager_id(ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_id),
    .io_network_acquire_ready(ClientTileLinkNetworkPort_1_io_network_acquire_ready),
    .io_network_acquire_valid(ClientTileLinkNetworkPort_1_io_network_acquire_valid),
    .io_network_acquire_bits_header_src(ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src),
    .io_network_acquire_bits_header_dst(ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst),
    .io_network_acquire_bits_payload_addr_block(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block),
    .io_network_acquire_bits_payload_client_xact_id(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id),
    .io_network_acquire_bits_payload_addr_beat(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat),
    .io_network_acquire_bits_payload_is_builtin_type(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type),
    .io_network_acquire_bits_payload_a_type(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type),
    .io_network_acquire_bits_payload_union(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union),
    .io_network_acquire_bits_payload_data(ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data),
    .io_network_grant_ready(ClientTileLinkNetworkPort_1_io_network_grant_ready),
    .io_network_grant_valid(ClientTileLinkNetworkPort_1_io_network_grant_valid),
    .io_network_grant_bits_header_src(ClientTileLinkNetworkPort_1_io_network_grant_bits_header_src),
    .io_network_grant_bits_header_dst(ClientTileLinkNetworkPort_1_io_network_grant_bits_header_dst),
    .io_network_grant_bits_payload_addr_beat(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat),
    .io_network_grant_bits_payload_client_xact_id(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id),
    .io_network_grant_bits_payload_manager_xact_id(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id),
    .io_network_grant_bits_payload_is_builtin_type(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type),
    .io_network_grant_bits_payload_g_type(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type),
    .io_network_grant_bits_payload_data(ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_data),
    .io_network_finish_ready(ClientTileLinkNetworkPort_1_io_network_finish_ready),
    .io_network_finish_valid(ClientTileLinkNetworkPort_1_io_network_finish_valid),
    .io_network_finish_bits_header_src(ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src),
    .io_network_finish_bits_header_dst(ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst),
    .io_network_finish_bits_payload_manager_xact_id(ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id),
    .io_network_probe_ready(ClientTileLinkNetworkPort_1_io_network_probe_ready),
    .io_network_probe_valid(ClientTileLinkNetworkPort_1_io_network_probe_valid),
    .io_network_probe_bits_header_src(ClientTileLinkNetworkPort_1_io_network_probe_bits_header_src),
    .io_network_probe_bits_header_dst(ClientTileLinkNetworkPort_1_io_network_probe_bits_header_dst),
    .io_network_probe_bits_payload_addr_block(ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block),
    .io_network_probe_bits_payload_p_type(ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type),
    .io_network_release_ready(ClientTileLinkNetworkPort_1_io_network_release_ready),
    .io_network_release_valid(ClientTileLinkNetworkPort_1_io_network_release_valid),
    .io_network_release_bits_header_src(ClientTileLinkNetworkPort_1_io_network_release_bits_header_src),
    .io_network_release_bits_header_dst(ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst),
    .io_network_release_bits_payload_addr_beat(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat),
    .io_network_release_bits_payload_addr_block(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block),
    .io_network_release_bits_payload_client_xact_id(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id),
    .io_network_release_bits_payload_voluntary(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary),
    .io_network_release_bits_payload_r_type(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type),
    .io_network_release_bits_payload_data(ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data)
  );
  TileLinkEnqueuer_1 TileLinkEnqueuer_1_1 (
    .clk(TileLinkEnqueuer_1_1_clk),
    .reset(TileLinkEnqueuer_1_1_reset),
    .io_client_acquire_ready(TileLinkEnqueuer_1_1_io_client_acquire_ready),
    .io_client_acquire_valid(TileLinkEnqueuer_1_1_io_client_acquire_valid),
    .io_client_acquire_bits_header_src(TileLinkEnqueuer_1_1_io_client_acquire_bits_header_src),
    .io_client_acquire_bits_header_dst(TileLinkEnqueuer_1_1_io_client_acquire_bits_header_dst),
    .io_client_acquire_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_block),
    .io_client_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_client_xact_id),
    .io_client_acquire_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_beat),
    .io_client_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_is_builtin_type),
    .io_client_acquire_bits_payload_a_type(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_a_type),
    .io_client_acquire_bits_payload_union(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_union),
    .io_client_acquire_bits_payload_data(TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_data),
    .io_client_grant_ready(TileLinkEnqueuer_1_1_io_client_grant_ready),
    .io_client_grant_valid(TileLinkEnqueuer_1_1_io_client_grant_valid),
    .io_client_grant_bits_header_src(TileLinkEnqueuer_1_1_io_client_grant_bits_header_src),
    .io_client_grant_bits_header_dst(TileLinkEnqueuer_1_1_io_client_grant_bits_header_dst),
    .io_client_grant_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_addr_beat),
    .io_client_grant_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_client_xact_id),
    .io_client_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_manager_xact_id),
    .io_client_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_is_builtin_type),
    .io_client_grant_bits_payload_g_type(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_g_type),
    .io_client_grant_bits_payload_data(TileLinkEnqueuer_1_1_io_client_grant_bits_payload_data),
    .io_client_finish_ready(TileLinkEnqueuer_1_1_io_client_finish_ready),
    .io_client_finish_valid(TileLinkEnqueuer_1_1_io_client_finish_valid),
    .io_client_finish_bits_header_src(TileLinkEnqueuer_1_1_io_client_finish_bits_header_src),
    .io_client_finish_bits_header_dst(TileLinkEnqueuer_1_1_io_client_finish_bits_header_dst),
    .io_client_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_1_1_io_client_finish_bits_payload_manager_xact_id),
    .io_client_probe_ready(TileLinkEnqueuer_1_1_io_client_probe_ready),
    .io_client_probe_valid(TileLinkEnqueuer_1_1_io_client_probe_valid),
    .io_client_probe_bits_header_src(TileLinkEnqueuer_1_1_io_client_probe_bits_header_src),
    .io_client_probe_bits_header_dst(TileLinkEnqueuer_1_1_io_client_probe_bits_header_dst),
    .io_client_probe_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_client_probe_bits_payload_addr_block),
    .io_client_probe_bits_payload_p_type(TileLinkEnqueuer_1_1_io_client_probe_bits_payload_p_type),
    .io_client_release_ready(TileLinkEnqueuer_1_1_io_client_release_ready),
    .io_client_release_valid(TileLinkEnqueuer_1_1_io_client_release_valid),
    .io_client_release_bits_header_src(TileLinkEnqueuer_1_1_io_client_release_bits_header_src),
    .io_client_release_bits_header_dst(TileLinkEnqueuer_1_1_io_client_release_bits_header_dst),
    .io_client_release_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_beat),
    .io_client_release_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_block),
    .io_client_release_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_client_release_bits_payload_client_xact_id),
    .io_client_release_bits_payload_voluntary(TileLinkEnqueuer_1_1_io_client_release_bits_payload_voluntary),
    .io_client_release_bits_payload_r_type(TileLinkEnqueuer_1_1_io_client_release_bits_payload_r_type),
    .io_client_release_bits_payload_data(TileLinkEnqueuer_1_1_io_client_release_bits_payload_data),
    .io_manager_acquire_ready(TileLinkEnqueuer_1_1_io_manager_acquire_ready),
    .io_manager_acquire_valid(TileLinkEnqueuer_1_1_io_manager_acquire_valid),
    .io_manager_acquire_bits_header_src(TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_src),
    .io_manager_acquire_bits_header_dst(TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_dst),
    .io_manager_acquire_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_block),
    .io_manager_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_client_xact_id),
    .io_manager_acquire_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_beat),
    .io_manager_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_is_builtin_type),
    .io_manager_acquire_bits_payload_a_type(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_a_type),
    .io_manager_acquire_bits_payload_union(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_union),
    .io_manager_acquire_bits_payload_data(TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_data),
    .io_manager_grant_ready(TileLinkEnqueuer_1_1_io_manager_grant_ready),
    .io_manager_grant_valid(TileLinkEnqueuer_1_1_io_manager_grant_valid),
    .io_manager_grant_bits_header_src(TileLinkEnqueuer_1_1_io_manager_grant_bits_header_src),
    .io_manager_grant_bits_header_dst(TileLinkEnqueuer_1_1_io_manager_grant_bits_header_dst),
    .io_manager_grant_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_addr_beat),
    .io_manager_grant_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_client_xact_id),
    .io_manager_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_manager_xact_id),
    .io_manager_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_is_builtin_type),
    .io_manager_grant_bits_payload_g_type(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_g_type),
    .io_manager_grant_bits_payload_data(TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_data),
    .io_manager_finish_ready(TileLinkEnqueuer_1_1_io_manager_finish_ready),
    .io_manager_finish_valid(TileLinkEnqueuer_1_1_io_manager_finish_valid),
    .io_manager_finish_bits_header_src(TileLinkEnqueuer_1_1_io_manager_finish_bits_header_src),
    .io_manager_finish_bits_header_dst(TileLinkEnqueuer_1_1_io_manager_finish_bits_header_dst),
    .io_manager_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_1_1_io_manager_finish_bits_payload_manager_xact_id),
    .io_manager_probe_ready(TileLinkEnqueuer_1_1_io_manager_probe_ready),
    .io_manager_probe_valid(TileLinkEnqueuer_1_1_io_manager_probe_valid),
    .io_manager_probe_bits_header_src(TileLinkEnqueuer_1_1_io_manager_probe_bits_header_src),
    .io_manager_probe_bits_header_dst(TileLinkEnqueuer_1_1_io_manager_probe_bits_header_dst),
    .io_manager_probe_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_addr_block),
    .io_manager_probe_bits_payload_p_type(TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_p_type),
    .io_manager_release_ready(TileLinkEnqueuer_1_1_io_manager_release_ready),
    .io_manager_release_valid(TileLinkEnqueuer_1_1_io_manager_release_valid),
    .io_manager_release_bits_header_src(TileLinkEnqueuer_1_1_io_manager_release_bits_header_src),
    .io_manager_release_bits_header_dst(TileLinkEnqueuer_1_1_io_manager_release_bits_header_dst),
    .io_manager_release_bits_payload_addr_beat(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_beat),
    .io_manager_release_bits_payload_addr_block(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_block),
    .io_manager_release_bits_payload_client_xact_id(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_client_xact_id),
    .io_manager_release_bits_payload_voluntary(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_voluntary),
    .io_manager_release_bits_payload_r_type(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_r_type),
    .io_manager_release_bits_payload_data(TileLinkEnqueuer_1_1_io_manager_release_bits_payload_data)
  );
  ClientUncachedTileLinkNetworkPort ClientUncachedTileLinkNetworkPort_1 (
    .clk(ClientUncachedTileLinkNetworkPort_1_clk),
    .reset(ClientUncachedTileLinkNetworkPort_1_reset),
    .io_client_acquire_ready(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_ready),
    .io_client_acquire_valid(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_valid),
    .io_client_acquire_bits_addr_block(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_block),
    .io_client_acquire_bits_client_xact_id(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id),
    .io_client_acquire_bits_addr_beat(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat),
    .io_client_acquire_bits_is_builtin_type(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type),
    .io_client_acquire_bits_a_type(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_a_type),
    .io_client_acquire_bits_union(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_union),
    .io_client_acquire_bits_data(ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_data),
    .io_client_grant_ready(ClientUncachedTileLinkNetworkPort_1_io_client_grant_ready),
    .io_client_grant_valid(ClientUncachedTileLinkNetworkPort_1_io_client_grant_valid),
    .io_client_grant_bits_addr_beat(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_addr_beat),
    .io_client_grant_bits_client_xact_id(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id),
    .io_client_grant_bits_manager_xact_id(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id),
    .io_client_grant_bits_is_builtin_type(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type),
    .io_client_grant_bits_g_type(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_g_type),
    .io_client_grant_bits_data(ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_data),
    .io_network_acquire_ready(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_ready),
    .io_network_acquire_valid(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_valid),
    .io_network_acquire_bits_header_src(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_src),
    .io_network_acquire_bits_header_dst(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_dst),
    .io_network_acquire_bits_payload_addr_block(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block),
    .io_network_acquire_bits_payload_client_xact_id(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id),
    .io_network_acquire_bits_payload_addr_beat(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat),
    .io_network_acquire_bits_payload_is_builtin_type(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type),
    .io_network_acquire_bits_payload_a_type(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type),
    .io_network_acquire_bits_payload_union(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_union),
    .io_network_acquire_bits_payload_data(ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_data),
    .io_network_grant_ready(ClientUncachedTileLinkNetworkPort_1_io_network_grant_ready),
    .io_network_grant_valid(ClientUncachedTileLinkNetworkPort_1_io_network_grant_valid),
    .io_network_grant_bits_header_src(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_src),
    .io_network_grant_bits_header_dst(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_dst),
    .io_network_grant_bits_payload_addr_beat(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat),
    .io_network_grant_bits_payload_client_xact_id(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id),
    .io_network_grant_bits_payload_manager_xact_id(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id),
    .io_network_grant_bits_payload_is_builtin_type(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type),
    .io_network_grant_bits_payload_g_type(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type),
    .io_network_grant_bits_payload_data(ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_data),
    .io_network_finish_ready(ClientUncachedTileLinkNetworkPort_1_io_network_finish_ready),
    .io_network_finish_valid(ClientUncachedTileLinkNetworkPort_1_io_network_finish_valid),
    .io_network_finish_bits_header_src(ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_src),
    .io_network_finish_bits_header_dst(ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_dst),
    .io_network_finish_bits_payload_manager_xact_id(ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id),
    .io_network_probe_ready(ClientUncachedTileLinkNetworkPort_1_io_network_probe_ready),
    .io_network_probe_valid(ClientUncachedTileLinkNetworkPort_1_io_network_probe_valid),
    .io_network_probe_bits_header_src(ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_src),
    .io_network_probe_bits_header_dst(ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_dst),
    .io_network_probe_bits_payload_addr_block(ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block),
    .io_network_probe_bits_payload_p_type(ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type),
    .io_network_release_ready(ClientUncachedTileLinkNetworkPort_1_io_network_release_ready),
    .io_network_release_valid(ClientUncachedTileLinkNetworkPort_1_io_network_release_valid),
    .io_network_release_bits_header_src(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_src),
    .io_network_release_bits_header_dst(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_dst),
    .io_network_release_bits_payload_addr_beat(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat),
    .io_network_release_bits_payload_addr_block(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block),
    .io_network_release_bits_payload_client_xact_id(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id),
    .io_network_release_bits_payload_voluntary(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary),
    .io_network_release_bits_payload_r_type(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_r_type),
    .io_network_release_bits_payload_data(ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_data)
  );
  ManagerTileLinkNetworkPort ManagerTileLinkNetworkPort_2 (
    .clk(ManagerTileLinkNetworkPort_2_clk),
    .reset(ManagerTileLinkNetworkPort_2_reset),
    .io_manager_acquire_ready(ManagerTileLinkNetworkPort_2_io_manager_acquire_ready),
    .io_manager_acquire_valid(ManagerTileLinkNetworkPort_2_io_manager_acquire_valid),
    .io_manager_acquire_bits_addr_block(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_block),
    .io_manager_acquire_bits_client_xact_id(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_xact_id),
    .io_manager_acquire_bits_addr_beat(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_beat),
    .io_manager_acquire_bits_is_builtin_type(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_is_builtin_type),
    .io_manager_acquire_bits_a_type(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_a_type),
    .io_manager_acquire_bits_union(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_union),
    .io_manager_acquire_bits_data(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_data),
    .io_manager_acquire_bits_client_id(ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_id),
    .io_manager_grant_ready(ManagerTileLinkNetworkPort_2_io_manager_grant_ready),
    .io_manager_grant_valid(ManagerTileLinkNetworkPort_2_io_manager_grant_valid),
    .io_manager_grant_bits_addr_beat(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_addr_beat),
    .io_manager_grant_bits_client_xact_id(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_xact_id),
    .io_manager_grant_bits_manager_xact_id(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_manager_xact_id),
    .io_manager_grant_bits_is_builtin_type(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_is_builtin_type),
    .io_manager_grant_bits_g_type(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_g_type),
    .io_manager_grant_bits_data(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_data),
    .io_manager_grant_bits_client_id(ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_id),
    .io_manager_finish_ready(ManagerTileLinkNetworkPort_2_io_manager_finish_ready),
    .io_manager_finish_valid(ManagerTileLinkNetworkPort_2_io_manager_finish_valid),
    .io_manager_finish_bits_manager_xact_id(ManagerTileLinkNetworkPort_2_io_manager_finish_bits_manager_xact_id),
    .io_manager_probe_ready(ManagerTileLinkNetworkPort_2_io_manager_probe_ready),
    .io_manager_probe_valid(ManagerTileLinkNetworkPort_2_io_manager_probe_valid),
    .io_manager_probe_bits_addr_block(ManagerTileLinkNetworkPort_2_io_manager_probe_bits_addr_block),
    .io_manager_probe_bits_p_type(ManagerTileLinkNetworkPort_2_io_manager_probe_bits_p_type),
    .io_manager_probe_bits_client_id(ManagerTileLinkNetworkPort_2_io_manager_probe_bits_client_id),
    .io_manager_release_ready(ManagerTileLinkNetworkPort_2_io_manager_release_ready),
    .io_manager_release_valid(ManagerTileLinkNetworkPort_2_io_manager_release_valid),
    .io_manager_release_bits_addr_beat(ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_beat),
    .io_manager_release_bits_addr_block(ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_block),
    .io_manager_release_bits_client_xact_id(ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_xact_id),
    .io_manager_release_bits_voluntary(ManagerTileLinkNetworkPort_2_io_manager_release_bits_voluntary),
    .io_manager_release_bits_r_type(ManagerTileLinkNetworkPort_2_io_manager_release_bits_r_type),
    .io_manager_release_bits_data(ManagerTileLinkNetworkPort_2_io_manager_release_bits_data),
    .io_manager_release_bits_client_id(ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_id),
    .io_network_acquire_ready(ManagerTileLinkNetworkPort_2_io_network_acquire_ready),
    .io_network_acquire_valid(ManagerTileLinkNetworkPort_2_io_network_acquire_valid),
    .io_network_acquire_bits_header_src(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_src),
    .io_network_acquire_bits_header_dst(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_dst),
    .io_network_acquire_bits_payload_addr_block(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block),
    .io_network_acquire_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id),
    .io_network_acquire_bits_payload_addr_beat(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat),
    .io_network_acquire_bits_payload_is_builtin_type(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type),
    .io_network_acquire_bits_payload_a_type(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type),
    .io_network_acquire_bits_payload_union(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_union),
    .io_network_acquire_bits_payload_data(ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_data),
    .io_network_grant_ready(ManagerTileLinkNetworkPort_2_io_network_grant_ready),
    .io_network_grant_valid(ManagerTileLinkNetworkPort_2_io_network_grant_valid),
    .io_network_grant_bits_header_src(ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_src),
    .io_network_grant_bits_header_dst(ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_dst),
    .io_network_grant_bits_payload_addr_beat(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_addr_beat),
    .io_network_grant_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_client_xact_id),
    .io_network_grant_bits_payload_manager_xact_id(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_manager_xact_id),
    .io_network_grant_bits_payload_is_builtin_type(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_is_builtin_type),
    .io_network_grant_bits_payload_g_type(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_g_type),
    .io_network_grant_bits_payload_data(ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_data),
    .io_network_finish_ready(ManagerTileLinkNetworkPort_2_io_network_finish_ready),
    .io_network_finish_valid(ManagerTileLinkNetworkPort_2_io_network_finish_valid),
    .io_network_finish_bits_header_src(ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_src),
    .io_network_finish_bits_header_dst(ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_dst),
    .io_network_finish_bits_payload_manager_xact_id(ManagerTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id),
    .io_network_probe_ready(ManagerTileLinkNetworkPort_2_io_network_probe_ready),
    .io_network_probe_valid(ManagerTileLinkNetworkPort_2_io_network_probe_valid),
    .io_network_probe_bits_header_src(ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_src),
    .io_network_probe_bits_header_dst(ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_dst),
    .io_network_probe_bits_payload_addr_block(ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_addr_block),
    .io_network_probe_bits_payload_p_type(ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_p_type),
    .io_network_release_ready(ManagerTileLinkNetworkPort_2_io_network_release_ready),
    .io_network_release_valid(ManagerTileLinkNetworkPort_2_io_network_release_valid),
    .io_network_release_bits_header_src(ManagerTileLinkNetworkPort_2_io_network_release_bits_header_src),
    .io_network_release_bits_header_dst(ManagerTileLinkNetworkPort_2_io_network_release_bits_header_dst),
    .io_network_release_bits_payload_addr_beat(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat),
    .io_network_release_bits_payload_addr_block(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block),
    .io_network_release_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id),
    .io_network_release_bits_payload_voluntary(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary),
    .io_network_release_bits_payload_r_type(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_r_type),
    .io_network_release_bits_payload_data(ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_data)
  );
  TileLinkEnqueuer_2 TileLinkEnqueuer_2_1 (
    .clk(TileLinkEnqueuer_2_1_clk),
    .reset(TileLinkEnqueuer_2_1_reset),
    .io_client_acquire_ready(TileLinkEnqueuer_2_1_io_client_acquire_ready),
    .io_client_acquire_valid(TileLinkEnqueuer_2_1_io_client_acquire_valid),
    .io_client_acquire_bits_header_src(TileLinkEnqueuer_2_1_io_client_acquire_bits_header_src),
    .io_client_acquire_bits_header_dst(TileLinkEnqueuer_2_1_io_client_acquire_bits_header_dst),
    .io_client_acquire_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_block),
    .io_client_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_client_xact_id),
    .io_client_acquire_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_beat),
    .io_client_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_is_builtin_type),
    .io_client_acquire_bits_payload_a_type(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_a_type),
    .io_client_acquire_bits_payload_union(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_union),
    .io_client_acquire_bits_payload_data(TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_data),
    .io_client_grant_ready(TileLinkEnqueuer_2_1_io_client_grant_ready),
    .io_client_grant_valid(TileLinkEnqueuer_2_1_io_client_grant_valid),
    .io_client_grant_bits_header_src(TileLinkEnqueuer_2_1_io_client_grant_bits_header_src),
    .io_client_grant_bits_header_dst(TileLinkEnqueuer_2_1_io_client_grant_bits_header_dst),
    .io_client_grant_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_addr_beat),
    .io_client_grant_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_client_xact_id),
    .io_client_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_manager_xact_id),
    .io_client_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_is_builtin_type),
    .io_client_grant_bits_payload_g_type(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_g_type),
    .io_client_grant_bits_payload_data(TileLinkEnqueuer_2_1_io_client_grant_bits_payload_data),
    .io_client_finish_ready(TileLinkEnqueuer_2_1_io_client_finish_ready),
    .io_client_finish_valid(TileLinkEnqueuer_2_1_io_client_finish_valid),
    .io_client_finish_bits_header_src(TileLinkEnqueuer_2_1_io_client_finish_bits_header_src),
    .io_client_finish_bits_header_dst(TileLinkEnqueuer_2_1_io_client_finish_bits_header_dst),
    .io_client_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_2_1_io_client_finish_bits_payload_manager_xact_id),
    .io_client_probe_ready(TileLinkEnqueuer_2_1_io_client_probe_ready),
    .io_client_probe_valid(TileLinkEnqueuer_2_1_io_client_probe_valid),
    .io_client_probe_bits_header_src(TileLinkEnqueuer_2_1_io_client_probe_bits_header_src),
    .io_client_probe_bits_header_dst(TileLinkEnqueuer_2_1_io_client_probe_bits_header_dst),
    .io_client_probe_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_client_probe_bits_payload_addr_block),
    .io_client_probe_bits_payload_p_type(TileLinkEnqueuer_2_1_io_client_probe_bits_payload_p_type),
    .io_client_release_ready(TileLinkEnqueuer_2_1_io_client_release_ready),
    .io_client_release_valid(TileLinkEnqueuer_2_1_io_client_release_valid),
    .io_client_release_bits_header_src(TileLinkEnqueuer_2_1_io_client_release_bits_header_src),
    .io_client_release_bits_header_dst(TileLinkEnqueuer_2_1_io_client_release_bits_header_dst),
    .io_client_release_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_beat),
    .io_client_release_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_block),
    .io_client_release_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_client_release_bits_payload_client_xact_id),
    .io_client_release_bits_payload_voluntary(TileLinkEnqueuer_2_1_io_client_release_bits_payload_voluntary),
    .io_client_release_bits_payload_r_type(TileLinkEnqueuer_2_1_io_client_release_bits_payload_r_type),
    .io_client_release_bits_payload_data(TileLinkEnqueuer_2_1_io_client_release_bits_payload_data),
    .io_manager_acquire_ready(TileLinkEnqueuer_2_1_io_manager_acquire_ready),
    .io_manager_acquire_valid(TileLinkEnqueuer_2_1_io_manager_acquire_valid),
    .io_manager_acquire_bits_header_src(TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_src),
    .io_manager_acquire_bits_header_dst(TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_dst),
    .io_manager_acquire_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_block),
    .io_manager_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_client_xact_id),
    .io_manager_acquire_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_beat),
    .io_manager_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_is_builtin_type),
    .io_manager_acquire_bits_payload_a_type(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_a_type),
    .io_manager_acquire_bits_payload_union(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_union),
    .io_manager_acquire_bits_payload_data(TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_data),
    .io_manager_grant_ready(TileLinkEnqueuer_2_1_io_manager_grant_ready),
    .io_manager_grant_valid(TileLinkEnqueuer_2_1_io_manager_grant_valid),
    .io_manager_grant_bits_header_src(TileLinkEnqueuer_2_1_io_manager_grant_bits_header_src),
    .io_manager_grant_bits_header_dst(TileLinkEnqueuer_2_1_io_manager_grant_bits_header_dst),
    .io_manager_grant_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_addr_beat),
    .io_manager_grant_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_client_xact_id),
    .io_manager_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_manager_xact_id),
    .io_manager_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_is_builtin_type),
    .io_manager_grant_bits_payload_g_type(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_g_type),
    .io_manager_grant_bits_payload_data(TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_data),
    .io_manager_finish_ready(TileLinkEnqueuer_2_1_io_manager_finish_ready),
    .io_manager_finish_valid(TileLinkEnqueuer_2_1_io_manager_finish_valid),
    .io_manager_finish_bits_header_src(TileLinkEnqueuer_2_1_io_manager_finish_bits_header_src),
    .io_manager_finish_bits_header_dst(TileLinkEnqueuer_2_1_io_manager_finish_bits_header_dst),
    .io_manager_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_2_1_io_manager_finish_bits_payload_manager_xact_id),
    .io_manager_probe_ready(TileLinkEnqueuer_2_1_io_manager_probe_ready),
    .io_manager_probe_valid(TileLinkEnqueuer_2_1_io_manager_probe_valid),
    .io_manager_probe_bits_header_src(TileLinkEnqueuer_2_1_io_manager_probe_bits_header_src),
    .io_manager_probe_bits_header_dst(TileLinkEnqueuer_2_1_io_manager_probe_bits_header_dst),
    .io_manager_probe_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_addr_block),
    .io_manager_probe_bits_payload_p_type(TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_p_type),
    .io_manager_release_ready(TileLinkEnqueuer_2_1_io_manager_release_ready),
    .io_manager_release_valid(TileLinkEnqueuer_2_1_io_manager_release_valid),
    .io_manager_release_bits_header_src(TileLinkEnqueuer_2_1_io_manager_release_bits_header_src),
    .io_manager_release_bits_header_dst(TileLinkEnqueuer_2_1_io_manager_release_bits_header_dst),
    .io_manager_release_bits_payload_addr_beat(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_beat),
    .io_manager_release_bits_payload_addr_block(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_block),
    .io_manager_release_bits_payload_client_xact_id(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_client_xact_id),
    .io_manager_release_bits_payload_voluntary(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_voluntary),
    .io_manager_release_bits_payload_r_type(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_r_type),
    .io_manager_release_bits_payload_data(TileLinkEnqueuer_2_1_io_manager_release_bits_payload_data)
  );
  ManagerTileLinkNetworkPort_1 ManagerTileLinkNetworkPort_1_1 (
    .clk(ManagerTileLinkNetworkPort_1_1_clk),
    .reset(ManagerTileLinkNetworkPort_1_1_reset),
    .io_manager_acquire_ready(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_ready),
    .io_manager_acquire_valid(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_valid),
    .io_manager_acquire_bits_addr_block(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_block),
    .io_manager_acquire_bits_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_xact_id),
    .io_manager_acquire_bits_addr_beat(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_beat),
    .io_manager_acquire_bits_is_builtin_type(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_is_builtin_type),
    .io_manager_acquire_bits_a_type(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_a_type),
    .io_manager_acquire_bits_union(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_union),
    .io_manager_acquire_bits_data(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_data),
    .io_manager_acquire_bits_client_id(ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_id),
    .io_manager_grant_ready(ManagerTileLinkNetworkPort_1_1_io_manager_grant_ready),
    .io_manager_grant_valid(ManagerTileLinkNetworkPort_1_1_io_manager_grant_valid),
    .io_manager_grant_bits_addr_beat(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_addr_beat),
    .io_manager_grant_bits_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_xact_id),
    .io_manager_grant_bits_manager_xact_id(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_manager_xact_id),
    .io_manager_grant_bits_is_builtin_type(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_is_builtin_type),
    .io_manager_grant_bits_g_type(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_g_type),
    .io_manager_grant_bits_data(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_data),
    .io_manager_grant_bits_client_id(ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_id),
    .io_manager_finish_ready(ManagerTileLinkNetworkPort_1_1_io_manager_finish_ready),
    .io_manager_finish_valid(ManagerTileLinkNetworkPort_1_1_io_manager_finish_valid),
    .io_manager_finish_bits_manager_xact_id(ManagerTileLinkNetworkPort_1_1_io_manager_finish_bits_manager_xact_id),
    .io_manager_probe_ready(ManagerTileLinkNetworkPort_1_1_io_manager_probe_ready),
    .io_manager_probe_valid(ManagerTileLinkNetworkPort_1_1_io_manager_probe_valid),
    .io_manager_probe_bits_addr_block(ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_addr_block),
    .io_manager_probe_bits_p_type(ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_p_type),
    .io_manager_probe_bits_client_id(ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_client_id),
    .io_manager_release_ready(ManagerTileLinkNetworkPort_1_1_io_manager_release_ready),
    .io_manager_release_valid(ManagerTileLinkNetworkPort_1_1_io_manager_release_valid),
    .io_manager_release_bits_addr_beat(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_beat),
    .io_manager_release_bits_addr_block(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_block),
    .io_manager_release_bits_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_xact_id),
    .io_manager_release_bits_voluntary(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_voluntary),
    .io_manager_release_bits_r_type(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_r_type),
    .io_manager_release_bits_data(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_data),
    .io_manager_release_bits_client_id(ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_id),
    .io_network_acquire_ready(ManagerTileLinkNetworkPort_1_1_io_network_acquire_ready),
    .io_network_acquire_valid(ManagerTileLinkNetworkPort_1_1_io_network_acquire_valid),
    .io_network_acquire_bits_header_src(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_src),
    .io_network_acquire_bits_header_dst(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_dst),
    .io_network_acquire_bits_payload_addr_block(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_block),
    .io_network_acquire_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_client_xact_id),
    .io_network_acquire_bits_payload_addr_beat(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_beat),
    .io_network_acquire_bits_payload_is_builtin_type(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_is_builtin_type),
    .io_network_acquire_bits_payload_a_type(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_a_type),
    .io_network_acquire_bits_payload_union(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_union),
    .io_network_acquire_bits_payload_data(ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_data),
    .io_network_grant_ready(ManagerTileLinkNetworkPort_1_1_io_network_grant_ready),
    .io_network_grant_valid(ManagerTileLinkNetworkPort_1_1_io_network_grant_valid),
    .io_network_grant_bits_header_src(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_src),
    .io_network_grant_bits_header_dst(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_dst),
    .io_network_grant_bits_payload_addr_beat(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_addr_beat),
    .io_network_grant_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_client_xact_id),
    .io_network_grant_bits_payload_manager_xact_id(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_manager_xact_id),
    .io_network_grant_bits_payload_is_builtin_type(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_is_builtin_type),
    .io_network_grant_bits_payload_g_type(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_g_type),
    .io_network_grant_bits_payload_data(ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_data),
    .io_network_finish_ready(ManagerTileLinkNetworkPort_1_1_io_network_finish_ready),
    .io_network_finish_valid(ManagerTileLinkNetworkPort_1_1_io_network_finish_valid),
    .io_network_finish_bits_header_src(ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_src),
    .io_network_finish_bits_header_dst(ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_dst),
    .io_network_finish_bits_payload_manager_xact_id(ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_payload_manager_xact_id),
    .io_network_probe_ready(ManagerTileLinkNetworkPort_1_1_io_network_probe_ready),
    .io_network_probe_valid(ManagerTileLinkNetworkPort_1_1_io_network_probe_valid),
    .io_network_probe_bits_header_src(ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_src),
    .io_network_probe_bits_header_dst(ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_dst),
    .io_network_probe_bits_payload_addr_block(ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_addr_block),
    .io_network_probe_bits_payload_p_type(ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_p_type),
    .io_network_release_ready(ManagerTileLinkNetworkPort_1_1_io_network_release_ready),
    .io_network_release_valid(ManagerTileLinkNetworkPort_1_1_io_network_release_valid),
    .io_network_release_bits_header_src(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_src),
    .io_network_release_bits_header_dst(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_dst),
    .io_network_release_bits_payload_addr_beat(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_beat),
    .io_network_release_bits_payload_addr_block(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_block),
    .io_network_release_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_client_xact_id),
    .io_network_release_bits_payload_voluntary(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_voluntary),
    .io_network_release_bits_payload_r_type(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_r_type),
    .io_network_release_bits_payload_data(ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_data)
  );
  TileLinkEnqueuer_2 TileLinkEnqueuer_3_1 (
    .clk(TileLinkEnqueuer_3_1_clk),
    .reset(TileLinkEnqueuer_3_1_reset),
    .io_client_acquire_ready(TileLinkEnqueuer_3_1_io_client_acquire_ready),
    .io_client_acquire_valid(TileLinkEnqueuer_3_1_io_client_acquire_valid),
    .io_client_acquire_bits_header_src(TileLinkEnqueuer_3_1_io_client_acquire_bits_header_src),
    .io_client_acquire_bits_header_dst(TileLinkEnqueuer_3_1_io_client_acquire_bits_header_dst),
    .io_client_acquire_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_block),
    .io_client_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_client_xact_id),
    .io_client_acquire_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_beat),
    .io_client_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_is_builtin_type),
    .io_client_acquire_bits_payload_a_type(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_a_type),
    .io_client_acquire_bits_payload_union(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_union),
    .io_client_acquire_bits_payload_data(TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_data),
    .io_client_grant_ready(TileLinkEnqueuer_3_1_io_client_grant_ready),
    .io_client_grant_valid(TileLinkEnqueuer_3_1_io_client_grant_valid),
    .io_client_grant_bits_header_src(TileLinkEnqueuer_3_1_io_client_grant_bits_header_src),
    .io_client_grant_bits_header_dst(TileLinkEnqueuer_3_1_io_client_grant_bits_header_dst),
    .io_client_grant_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_addr_beat),
    .io_client_grant_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_client_xact_id),
    .io_client_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_manager_xact_id),
    .io_client_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_is_builtin_type),
    .io_client_grant_bits_payload_g_type(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_g_type),
    .io_client_grant_bits_payload_data(TileLinkEnqueuer_3_1_io_client_grant_bits_payload_data),
    .io_client_finish_ready(TileLinkEnqueuer_3_1_io_client_finish_ready),
    .io_client_finish_valid(TileLinkEnqueuer_3_1_io_client_finish_valid),
    .io_client_finish_bits_header_src(TileLinkEnqueuer_3_1_io_client_finish_bits_header_src),
    .io_client_finish_bits_header_dst(TileLinkEnqueuer_3_1_io_client_finish_bits_header_dst),
    .io_client_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_3_1_io_client_finish_bits_payload_manager_xact_id),
    .io_client_probe_ready(TileLinkEnqueuer_3_1_io_client_probe_ready),
    .io_client_probe_valid(TileLinkEnqueuer_3_1_io_client_probe_valid),
    .io_client_probe_bits_header_src(TileLinkEnqueuer_3_1_io_client_probe_bits_header_src),
    .io_client_probe_bits_header_dst(TileLinkEnqueuer_3_1_io_client_probe_bits_header_dst),
    .io_client_probe_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_client_probe_bits_payload_addr_block),
    .io_client_probe_bits_payload_p_type(TileLinkEnqueuer_3_1_io_client_probe_bits_payload_p_type),
    .io_client_release_ready(TileLinkEnqueuer_3_1_io_client_release_ready),
    .io_client_release_valid(TileLinkEnqueuer_3_1_io_client_release_valid),
    .io_client_release_bits_header_src(TileLinkEnqueuer_3_1_io_client_release_bits_header_src),
    .io_client_release_bits_header_dst(TileLinkEnqueuer_3_1_io_client_release_bits_header_dst),
    .io_client_release_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_beat),
    .io_client_release_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_block),
    .io_client_release_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_client_release_bits_payload_client_xact_id),
    .io_client_release_bits_payload_voluntary(TileLinkEnqueuer_3_1_io_client_release_bits_payload_voluntary),
    .io_client_release_bits_payload_r_type(TileLinkEnqueuer_3_1_io_client_release_bits_payload_r_type),
    .io_client_release_bits_payload_data(TileLinkEnqueuer_3_1_io_client_release_bits_payload_data),
    .io_manager_acquire_ready(TileLinkEnqueuer_3_1_io_manager_acquire_ready),
    .io_manager_acquire_valid(TileLinkEnqueuer_3_1_io_manager_acquire_valid),
    .io_manager_acquire_bits_header_src(TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_src),
    .io_manager_acquire_bits_header_dst(TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_dst),
    .io_manager_acquire_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_block),
    .io_manager_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_client_xact_id),
    .io_manager_acquire_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_beat),
    .io_manager_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_is_builtin_type),
    .io_manager_acquire_bits_payload_a_type(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_a_type),
    .io_manager_acquire_bits_payload_union(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_union),
    .io_manager_acquire_bits_payload_data(TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_data),
    .io_manager_grant_ready(TileLinkEnqueuer_3_1_io_manager_grant_ready),
    .io_manager_grant_valid(TileLinkEnqueuer_3_1_io_manager_grant_valid),
    .io_manager_grant_bits_header_src(TileLinkEnqueuer_3_1_io_manager_grant_bits_header_src),
    .io_manager_grant_bits_header_dst(TileLinkEnqueuer_3_1_io_manager_grant_bits_header_dst),
    .io_manager_grant_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_addr_beat),
    .io_manager_grant_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_client_xact_id),
    .io_manager_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_manager_xact_id),
    .io_manager_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_is_builtin_type),
    .io_manager_grant_bits_payload_g_type(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_g_type),
    .io_manager_grant_bits_payload_data(TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_data),
    .io_manager_finish_ready(TileLinkEnqueuer_3_1_io_manager_finish_ready),
    .io_manager_finish_valid(TileLinkEnqueuer_3_1_io_manager_finish_valid),
    .io_manager_finish_bits_header_src(TileLinkEnqueuer_3_1_io_manager_finish_bits_header_src),
    .io_manager_finish_bits_header_dst(TileLinkEnqueuer_3_1_io_manager_finish_bits_header_dst),
    .io_manager_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_3_1_io_manager_finish_bits_payload_manager_xact_id),
    .io_manager_probe_ready(TileLinkEnqueuer_3_1_io_manager_probe_ready),
    .io_manager_probe_valid(TileLinkEnqueuer_3_1_io_manager_probe_valid),
    .io_manager_probe_bits_header_src(TileLinkEnqueuer_3_1_io_manager_probe_bits_header_src),
    .io_manager_probe_bits_header_dst(TileLinkEnqueuer_3_1_io_manager_probe_bits_header_dst),
    .io_manager_probe_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_addr_block),
    .io_manager_probe_bits_payload_p_type(TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_p_type),
    .io_manager_release_ready(TileLinkEnqueuer_3_1_io_manager_release_ready),
    .io_manager_release_valid(TileLinkEnqueuer_3_1_io_manager_release_valid),
    .io_manager_release_bits_header_src(TileLinkEnqueuer_3_1_io_manager_release_bits_header_src),
    .io_manager_release_bits_header_dst(TileLinkEnqueuer_3_1_io_manager_release_bits_header_dst),
    .io_manager_release_bits_payload_addr_beat(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_beat),
    .io_manager_release_bits_payload_addr_block(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_block),
    .io_manager_release_bits_payload_client_xact_id(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_client_xact_id),
    .io_manager_release_bits_payload_voluntary(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_voluntary),
    .io_manager_release_bits_payload_r_type(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_r_type),
    .io_manager_release_bits_payload_data(TileLinkEnqueuer_3_1_io_manager_release_bits_payload_data)
  );
  BasicBus acqNet (
    .clk(acqNet_clk),
    .reset(acqNet_reset),
    .io_in_0_ready(acqNet_io_in_0_ready),
    .io_in_0_valid(acqNet_io_in_0_valid),
    .io_in_0_bits_header_src(acqNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(acqNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_block(acqNet_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_client_xact_id(acqNet_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_addr_beat(acqNet_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_is_builtin_type(acqNet_io_in_0_bits_payload_is_builtin_type),
    .io_in_0_bits_payload_a_type(acqNet_io_in_0_bits_payload_a_type),
    .io_in_0_bits_payload_union(acqNet_io_in_0_bits_payload_union),
    .io_in_0_bits_payload_data(acqNet_io_in_0_bits_payload_data),
    .io_in_1_ready(acqNet_io_in_1_ready),
    .io_in_1_valid(acqNet_io_in_1_valid),
    .io_in_1_bits_header_src(acqNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(acqNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_block(acqNet_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_client_xact_id(acqNet_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_addr_beat(acqNet_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_is_builtin_type(acqNet_io_in_1_bits_payload_is_builtin_type),
    .io_in_1_bits_payload_a_type(acqNet_io_in_1_bits_payload_a_type),
    .io_in_1_bits_payload_union(acqNet_io_in_1_bits_payload_union),
    .io_in_1_bits_payload_data(acqNet_io_in_1_bits_payload_data),
    .io_in_2_ready(acqNet_io_in_2_ready),
    .io_in_2_valid(acqNet_io_in_2_valid),
    .io_in_2_bits_header_src(acqNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(acqNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_block(acqNet_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_client_xact_id(acqNet_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_addr_beat(acqNet_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_is_builtin_type(acqNet_io_in_2_bits_payload_is_builtin_type),
    .io_in_2_bits_payload_a_type(acqNet_io_in_2_bits_payload_a_type),
    .io_in_2_bits_payload_union(acqNet_io_in_2_bits_payload_union),
    .io_in_2_bits_payload_data(acqNet_io_in_2_bits_payload_data),
    .io_in_3_ready(acqNet_io_in_3_ready),
    .io_in_3_valid(acqNet_io_in_3_valid),
    .io_in_3_bits_header_src(acqNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(acqNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_block(acqNet_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_client_xact_id(acqNet_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_addr_beat(acqNet_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_is_builtin_type(acqNet_io_in_3_bits_payload_is_builtin_type),
    .io_in_3_bits_payload_a_type(acqNet_io_in_3_bits_payload_a_type),
    .io_in_3_bits_payload_union(acqNet_io_in_3_bits_payload_union),
    .io_in_3_bits_payload_data(acqNet_io_in_3_bits_payload_data),
    .io_out_0_ready(acqNet_io_out_0_ready),
    .io_out_0_valid(acqNet_io_out_0_valid),
    .io_out_0_bits_header_src(acqNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(acqNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_addr_block(acqNet_io_out_0_bits_payload_addr_block),
    .io_out_0_bits_payload_client_xact_id(acqNet_io_out_0_bits_payload_client_xact_id),
    .io_out_0_bits_payload_addr_beat(acqNet_io_out_0_bits_payload_addr_beat),
    .io_out_0_bits_payload_is_builtin_type(acqNet_io_out_0_bits_payload_is_builtin_type),
    .io_out_0_bits_payload_a_type(acqNet_io_out_0_bits_payload_a_type),
    .io_out_0_bits_payload_union(acqNet_io_out_0_bits_payload_union),
    .io_out_0_bits_payload_data(acqNet_io_out_0_bits_payload_data),
    .io_out_1_ready(acqNet_io_out_1_ready),
    .io_out_1_valid(acqNet_io_out_1_valid),
    .io_out_1_bits_header_src(acqNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(acqNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_addr_block(acqNet_io_out_1_bits_payload_addr_block),
    .io_out_1_bits_payload_client_xact_id(acqNet_io_out_1_bits_payload_client_xact_id),
    .io_out_1_bits_payload_addr_beat(acqNet_io_out_1_bits_payload_addr_beat),
    .io_out_1_bits_payload_is_builtin_type(acqNet_io_out_1_bits_payload_is_builtin_type),
    .io_out_1_bits_payload_a_type(acqNet_io_out_1_bits_payload_a_type),
    .io_out_1_bits_payload_union(acqNet_io_out_1_bits_payload_union),
    .io_out_1_bits_payload_data(acqNet_io_out_1_bits_payload_data),
    .io_out_2_ready(acqNet_io_out_2_ready),
    .io_out_2_valid(acqNet_io_out_2_valid),
    .io_out_2_bits_header_src(acqNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(acqNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_addr_block(acqNet_io_out_2_bits_payload_addr_block),
    .io_out_2_bits_payload_client_xact_id(acqNet_io_out_2_bits_payload_client_xact_id),
    .io_out_2_bits_payload_addr_beat(acqNet_io_out_2_bits_payload_addr_beat),
    .io_out_2_bits_payload_is_builtin_type(acqNet_io_out_2_bits_payload_is_builtin_type),
    .io_out_2_bits_payload_a_type(acqNet_io_out_2_bits_payload_a_type),
    .io_out_2_bits_payload_union(acqNet_io_out_2_bits_payload_union),
    .io_out_2_bits_payload_data(acqNet_io_out_2_bits_payload_data),
    .io_out_3_ready(acqNet_io_out_3_ready),
    .io_out_3_valid(acqNet_io_out_3_valid),
    .io_out_3_bits_header_src(acqNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(acqNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_addr_block(acqNet_io_out_3_bits_payload_addr_block),
    .io_out_3_bits_payload_client_xact_id(acqNet_io_out_3_bits_payload_client_xact_id),
    .io_out_3_bits_payload_addr_beat(acqNet_io_out_3_bits_payload_addr_beat),
    .io_out_3_bits_payload_is_builtin_type(acqNet_io_out_3_bits_payload_is_builtin_type),
    .io_out_3_bits_payload_a_type(acqNet_io_out_3_bits_payload_a_type),
    .io_out_3_bits_payload_union(acqNet_io_out_3_bits_payload_union),
    .io_out_3_bits_payload_data(acqNet_io_out_3_bits_payload_data)
  );
  BasicBus_1 relNet (
    .clk(relNet_clk),
    .reset(relNet_reset),
    .io_in_0_ready(relNet_io_in_0_ready),
    .io_in_0_valid(relNet_io_in_0_valid),
    .io_in_0_bits_header_src(relNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(relNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_beat(relNet_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_addr_block(relNet_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_client_xact_id(relNet_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_voluntary(relNet_io_in_0_bits_payload_voluntary),
    .io_in_0_bits_payload_r_type(relNet_io_in_0_bits_payload_r_type),
    .io_in_0_bits_payload_data(relNet_io_in_0_bits_payload_data),
    .io_in_1_ready(relNet_io_in_1_ready),
    .io_in_1_valid(relNet_io_in_1_valid),
    .io_in_1_bits_header_src(relNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(relNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_beat(relNet_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_addr_block(relNet_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_client_xact_id(relNet_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_voluntary(relNet_io_in_1_bits_payload_voluntary),
    .io_in_1_bits_payload_r_type(relNet_io_in_1_bits_payload_r_type),
    .io_in_1_bits_payload_data(relNet_io_in_1_bits_payload_data),
    .io_in_2_ready(relNet_io_in_2_ready),
    .io_in_2_valid(relNet_io_in_2_valid),
    .io_in_2_bits_header_src(relNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(relNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_beat(relNet_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_addr_block(relNet_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_client_xact_id(relNet_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_voluntary(relNet_io_in_2_bits_payload_voluntary),
    .io_in_2_bits_payload_r_type(relNet_io_in_2_bits_payload_r_type),
    .io_in_2_bits_payload_data(relNet_io_in_2_bits_payload_data),
    .io_in_3_ready(relNet_io_in_3_ready),
    .io_in_3_valid(relNet_io_in_3_valid),
    .io_in_3_bits_header_src(relNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(relNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_beat(relNet_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_addr_block(relNet_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_client_xact_id(relNet_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_voluntary(relNet_io_in_3_bits_payload_voluntary),
    .io_in_3_bits_payload_r_type(relNet_io_in_3_bits_payload_r_type),
    .io_in_3_bits_payload_data(relNet_io_in_3_bits_payload_data),
    .io_out_0_ready(relNet_io_out_0_ready),
    .io_out_0_valid(relNet_io_out_0_valid),
    .io_out_0_bits_header_src(relNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(relNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_addr_beat(relNet_io_out_0_bits_payload_addr_beat),
    .io_out_0_bits_payload_addr_block(relNet_io_out_0_bits_payload_addr_block),
    .io_out_0_bits_payload_client_xact_id(relNet_io_out_0_bits_payload_client_xact_id),
    .io_out_0_bits_payload_voluntary(relNet_io_out_0_bits_payload_voluntary),
    .io_out_0_bits_payload_r_type(relNet_io_out_0_bits_payload_r_type),
    .io_out_0_bits_payload_data(relNet_io_out_0_bits_payload_data),
    .io_out_1_ready(relNet_io_out_1_ready),
    .io_out_1_valid(relNet_io_out_1_valid),
    .io_out_1_bits_header_src(relNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(relNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_addr_beat(relNet_io_out_1_bits_payload_addr_beat),
    .io_out_1_bits_payload_addr_block(relNet_io_out_1_bits_payload_addr_block),
    .io_out_1_bits_payload_client_xact_id(relNet_io_out_1_bits_payload_client_xact_id),
    .io_out_1_bits_payload_voluntary(relNet_io_out_1_bits_payload_voluntary),
    .io_out_1_bits_payload_r_type(relNet_io_out_1_bits_payload_r_type),
    .io_out_1_bits_payload_data(relNet_io_out_1_bits_payload_data),
    .io_out_2_ready(relNet_io_out_2_ready),
    .io_out_2_valid(relNet_io_out_2_valid),
    .io_out_2_bits_header_src(relNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(relNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_addr_beat(relNet_io_out_2_bits_payload_addr_beat),
    .io_out_2_bits_payload_addr_block(relNet_io_out_2_bits_payload_addr_block),
    .io_out_2_bits_payload_client_xact_id(relNet_io_out_2_bits_payload_client_xact_id),
    .io_out_2_bits_payload_voluntary(relNet_io_out_2_bits_payload_voluntary),
    .io_out_2_bits_payload_r_type(relNet_io_out_2_bits_payload_r_type),
    .io_out_2_bits_payload_data(relNet_io_out_2_bits_payload_data),
    .io_out_3_ready(relNet_io_out_3_ready),
    .io_out_3_valid(relNet_io_out_3_valid),
    .io_out_3_bits_header_src(relNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(relNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_addr_beat(relNet_io_out_3_bits_payload_addr_beat),
    .io_out_3_bits_payload_addr_block(relNet_io_out_3_bits_payload_addr_block),
    .io_out_3_bits_payload_client_xact_id(relNet_io_out_3_bits_payload_client_xact_id),
    .io_out_3_bits_payload_voluntary(relNet_io_out_3_bits_payload_voluntary),
    .io_out_3_bits_payload_r_type(relNet_io_out_3_bits_payload_r_type),
    .io_out_3_bits_payload_data(relNet_io_out_3_bits_payload_data)
  );
  BasicBus_2 prbNet (
    .clk(prbNet_clk),
    .reset(prbNet_reset),
    .io_in_0_ready(prbNet_io_in_0_ready),
    .io_in_0_valid(prbNet_io_in_0_valid),
    .io_in_0_bits_header_src(prbNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(prbNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_block(prbNet_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_p_type(prbNet_io_in_0_bits_payload_p_type),
    .io_in_1_ready(prbNet_io_in_1_ready),
    .io_in_1_valid(prbNet_io_in_1_valid),
    .io_in_1_bits_header_src(prbNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(prbNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_block(prbNet_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_p_type(prbNet_io_in_1_bits_payload_p_type),
    .io_in_2_ready(prbNet_io_in_2_ready),
    .io_in_2_valid(prbNet_io_in_2_valid),
    .io_in_2_bits_header_src(prbNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(prbNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_block(prbNet_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_p_type(prbNet_io_in_2_bits_payload_p_type),
    .io_in_3_ready(prbNet_io_in_3_ready),
    .io_in_3_valid(prbNet_io_in_3_valid),
    .io_in_3_bits_header_src(prbNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(prbNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_block(prbNet_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_p_type(prbNet_io_in_3_bits_payload_p_type),
    .io_out_0_ready(prbNet_io_out_0_ready),
    .io_out_0_valid(prbNet_io_out_0_valid),
    .io_out_0_bits_header_src(prbNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(prbNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_addr_block(prbNet_io_out_0_bits_payload_addr_block),
    .io_out_0_bits_payload_p_type(prbNet_io_out_0_bits_payload_p_type),
    .io_out_1_ready(prbNet_io_out_1_ready),
    .io_out_1_valid(prbNet_io_out_1_valid),
    .io_out_1_bits_header_src(prbNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(prbNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_addr_block(prbNet_io_out_1_bits_payload_addr_block),
    .io_out_1_bits_payload_p_type(prbNet_io_out_1_bits_payload_p_type),
    .io_out_2_ready(prbNet_io_out_2_ready),
    .io_out_2_valid(prbNet_io_out_2_valid),
    .io_out_2_bits_header_src(prbNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(prbNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_addr_block(prbNet_io_out_2_bits_payload_addr_block),
    .io_out_2_bits_payload_p_type(prbNet_io_out_2_bits_payload_p_type),
    .io_out_3_ready(prbNet_io_out_3_ready),
    .io_out_3_valid(prbNet_io_out_3_valid),
    .io_out_3_bits_header_src(prbNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(prbNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_addr_block(prbNet_io_out_3_bits_payload_addr_block),
    .io_out_3_bits_payload_p_type(prbNet_io_out_3_bits_payload_p_type)
  );
  BasicBus_3 gntNet (
    .clk(gntNet_clk),
    .reset(gntNet_reset),
    .io_in_0_ready(gntNet_io_in_0_ready),
    .io_in_0_valid(gntNet_io_in_0_valid),
    .io_in_0_bits_header_src(gntNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(gntNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_beat(gntNet_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_client_xact_id(gntNet_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_manager_xact_id(gntNet_io_in_0_bits_payload_manager_xact_id),
    .io_in_0_bits_payload_is_builtin_type(gntNet_io_in_0_bits_payload_is_builtin_type),
    .io_in_0_bits_payload_g_type(gntNet_io_in_0_bits_payload_g_type),
    .io_in_0_bits_payload_data(gntNet_io_in_0_bits_payload_data),
    .io_in_1_ready(gntNet_io_in_1_ready),
    .io_in_1_valid(gntNet_io_in_1_valid),
    .io_in_1_bits_header_src(gntNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(gntNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_beat(gntNet_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_client_xact_id(gntNet_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_manager_xact_id(gntNet_io_in_1_bits_payload_manager_xact_id),
    .io_in_1_bits_payload_is_builtin_type(gntNet_io_in_1_bits_payload_is_builtin_type),
    .io_in_1_bits_payload_g_type(gntNet_io_in_1_bits_payload_g_type),
    .io_in_1_bits_payload_data(gntNet_io_in_1_bits_payload_data),
    .io_in_2_ready(gntNet_io_in_2_ready),
    .io_in_2_valid(gntNet_io_in_2_valid),
    .io_in_2_bits_header_src(gntNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(gntNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_beat(gntNet_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_client_xact_id(gntNet_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_manager_xact_id(gntNet_io_in_2_bits_payload_manager_xact_id),
    .io_in_2_bits_payload_is_builtin_type(gntNet_io_in_2_bits_payload_is_builtin_type),
    .io_in_2_bits_payload_g_type(gntNet_io_in_2_bits_payload_g_type),
    .io_in_2_bits_payload_data(gntNet_io_in_2_bits_payload_data),
    .io_in_3_ready(gntNet_io_in_3_ready),
    .io_in_3_valid(gntNet_io_in_3_valid),
    .io_in_3_bits_header_src(gntNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(gntNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_beat(gntNet_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_client_xact_id(gntNet_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_manager_xact_id(gntNet_io_in_3_bits_payload_manager_xact_id),
    .io_in_3_bits_payload_is_builtin_type(gntNet_io_in_3_bits_payload_is_builtin_type),
    .io_in_3_bits_payload_g_type(gntNet_io_in_3_bits_payload_g_type),
    .io_in_3_bits_payload_data(gntNet_io_in_3_bits_payload_data),
    .io_out_0_ready(gntNet_io_out_0_ready),
    .io_out_0_valid(gntNet_io_out_0_valid),
    .io_out_0_bits_header_src(gntNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(gntNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_addr_beat(gntNet_io_out_0_bits_payload_addr_beat),
    .io_out_0_bits_payload_client_xact_id(gntNet_io_out_0_bits_payload_client_xact_id),
    .io_out_0_bits_payload_manager_xact_id(gntNet_io_out_0_bits_payload_manager_xact_id),
    .io_out_0_bits_payload_is_builtin_type(gntNet_io_out_0_bits_payload_is_builtin_type),
    .io_out_0_bits_payload_g_type(gntNet_io_out_0_bits_payload_g_type),
    .io_out_0_bits_payload_data(gntNet_io_out_0_bits_payload_data),
    .io_out_1_ready(gntNet_io_out_1_ready),
    .io_out_1_valid(gntNet_io_out_1_valid),
    .io_out_1_bits_header_src(gntNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(gntNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_addr_beat(gntNet_io_out_1_bits_payload_addr_beat),
    .io_out_1_bits_payload_client_xact_id(gntNet_io_out_1_bits_payload_client_xact_id),
    .io_out_1_bits_payload_manager_xact_id(gntNet_io_out_1_bits_payload_manager_xact_id),
    .io_out_1_bits_payload_is_builtin_type(gntNet_io_out_1_bits_payload_is_builtin_type),
    .io_out_1_bits_payload_g_type(gntNet_io_out_1_bits_payload_g_type),
    .io_out_1_bits_payload_data(gntNet_io_out_1_bits_payload_data),
    .io_out_2_ready(gntNet_io_out_2_ready),
    .io_out_2_valid(gntNet_io_out_2_valid),
    .io_out_2_bits_header_src(gntNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(gntNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_addr_beat(gntNet_io_out_2_bits_payload_addr_beat),
    .io_out_2_bits_payload_client_xact_id(gntNet_io_out_2_bits_payload_client_xact_id),
    .io_out_2_bits_payload_manager_xact_id(gntNet_io_out_2_bits_payload_manager_xact_id),
    .io_out_2_bits_payload_is_builtin_type(gntNet_io_out_2_bits_payload_is_builtin_type),
    .io_out_2_bits_payload_g_type(gntNet_io_out_2_bits_payload_g_type),
    .io_out_2_bits_payload_data(gntNet_io_out_2_bits_payload_data),
    .io_out_3_ready(gntNet_io_out_3_ready),
    .io_out_3_valid(gntNet_io_out_3_valid),
    .io_out_3_bits_header_src(gntNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(gntNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_addr_beat(gntNet_io_out_3_bits_payload_addr_beat),
    .io_out_3_bits_payload_client_xact_id(gntNet_io_out_3_bits_payload_client_xact_id),
    .io_out_3_bits_payload_manager_xact_id(gntNet_io_out_3_bits_payload_manager_xact_id),
    .io_out_3_bits_payload_is_builtin_type(gntNet_io_out_3_bits_payload_is_builtin_type),
    .io_out_3_bits_payload_g_type(gntNet_io_out_3_bits_payload_g_type),
    .io_out_3_bits_payload_data(gntNet_io_out_3_bits_payload_data)
  );
  BasicBus_4 ackNet (
    .clk(ackNet_clk),
    .reset(ackNet_reset),
    .io_in_0_ready(ackNet_io_in_0_ready),
    .io_in_0_valid(ackNet_io_in_0_valid),
    .io_in_0_bits_header_src(ackNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(ackNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_manager_xact_id(ackNet_io_in_0_bits_payload_manager_xact_id),
    .io_in_1_ready(ackNet_io_in_1_ready),
    .io_in_1_valid(ackNet_io_in_1_valid),
    .io_in_1_bits_header_src(ackNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(ackNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_manager_xact_id(ackNet_io_in_1_bits_payload_manager_xact_id),
    .io_in_2_ready(ackNet_io_in_2_ready),
    .io_in_2_valid(ackNet_io_in_2_valid),
    .io_in_2_bits_header_src(ackNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(ackNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_manager_xact_id(ackNet_io_in_2_bits_payload_manager_xact_id),
    .io_in_3_ready(ackNet_io_in_3_ready),
    .io_in_3_valid(ackNet_io_in_3_valid),
    .io_in_3_bits_header_src(ackNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(ackNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_manager_xact_id(ackNet_io_in_3_bits_payload_manager_xact_id),
    .io_out_0_ready(ackNet_io_out_0_ready),
    .io_out_0_valid(ackNet_io_out_0_valid),
    .io_out_0_bits_header_src(ackNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(ackNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_manager_xact_id(ackNet_io_out_0_bits_payload_manager_xact_id),
    .io_out_1_ready(ackNet_io_out_1_ready),
    .io_out_1_valid(ackNet_io_out_1_valid),
    .io_out_1_bits_header_src(ackNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(ackNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_manager_xact_id(ackNet_io_out_1_bits_payload_manager_xact_id),
    .io_out_2_ready(ackNet_io_out_2_ready),
    .io_out_2_valid(ackNet_io_out_2_valid),
    .io_out_2_bits_header_src(ackNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(ackNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_manager_xact_id(ackNet_io_out_2_bits_payload_manager_xact_id),
    .io_out_3_ready(ackNet_io_out_3_ready),
    .io_out_3_valid(ackNet_io_out_3_valid),
    .io_out_3_bits_header_src(ackNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(ackNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_manager_xact_id(ackNet_io_out_3_bits_payload_manager_xact_id)
  );
  assign io_clients_cached_0_acquire_ready = ClientTileLinkNetworkPort_1_io_client_acquire_ready;
  assign io_clients_cached_0_probe_valid = ClientTileLinkNetworkPort_1_io_client_probe_valid;
  assign io_clients_cached_0_probe_bits_addr_block = ClientTileLinkNetworkPort_1_io_client_probe_bits_addr_block;
  assign io_clients_cached_0_probe_bits_p_type = ClientTileLinkNetworkPort_1_io_client_probe_bits_p_type;
  assign io_clients_cached_0_release_ready = ClientTileLinkNetworkPort_1_io_client_release_ready;
  assign io_clients_cached_0_grant_valid = ClientTileLinkNetworkPort_1_io_client_grant_valid;
  assign io_clients_cached_0_grant_bits_addr_beat = ClientTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  assign io_clients_cached_0_grant_bits_client_xact_id = ClientTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  assign io_clients_cached_0_grant_bits_manager_xact_id = ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  assign io_clients_cached_0_grant_bits_is_builtin_type = ClientTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  assign io_clients_cached_0_grant_bits_g_type = ClientTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  assign io_clients_cached_0_grant_bits_data = ClientTileLinkNetworkPort_1_io_client_grant_bits_data;
  assign io_clients_cached_0_grant_bits_manager_id = ClientTileLinkNetworkPort_1_io_client_grant_bits_manager_id;
  assign io_clients_cached_0_finish_ready = ClientTileLinkNetworkPort_1_io_client_finish_ready;
  assign io_clients_uncached_0_acquire_ready = ClientUncachedTileLinkNetworkPort_1_io_client_acquire_ready;
  assign io_clients_uncached_0_grant_valid = ClientUncachedTileLinkNetworkPort_1_io_client_grant_valid;
  assign io_clients_uncached_0_grant_bits_addr_beat = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_addr_beat;
  assign io_clients_uncached_0_grant_bits_client_xact_id = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_client_xact_id;
  assign io_clients_uncached_0_grant_bits_manager_xact_id = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_manager_xact_id;
  assign io_clients_uncached_0_grant_bits_is_builtin_type = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_is_builtin_type;
  assign io_clients_uncached_0_grant_bits_g_type = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_g_type;
  assign io_clients_uncached_0_grant_bits_data = ClientUncachedTileLinkNetworkPort_1_io_client_grant_bits_data;
  assign io_managers_0_acquire_valid = ManagerTileLinkNetworkPort_2_io_manager_acquire_valid;
  assign io_managers_0_acquire_bits_addr_block = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_block;
  assign io_managers_0_acquire_bits_client_xact_id = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_xact_id;
  assign io_managers_0_acquire_bits_addr_beat = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_addr_beat;
  assign io_managers_0_acquire_bits_is_builtin_type = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_is_builtin_type;
  assign io_managers_0_acquire_bits_a_type = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_a_type;
  assign io_managers_0_acquire_bits_union = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_union;
  assign io_managers_0_acquire_bits_data = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_data;
  assign io_managers_0_acquire_bits_client_id = ManagerTileLinkNetworkPort_2_io_manager_acquire_bits_client_id;
  assign io_managers_0_grant_ready = ManagerTileLinkNetworkPort_2_io_manager_grant_ready;
  assign io_managers_0_finish_valid = ManagerTileLinkNetworkPort_2_io_manager_finish_valid;
  assign io_managers_0_finish_bits_manager_xact_id = ManagerTileLinkNetworkPort_2_io_manager_finish_bits_manager_xact_id;
  assign io_managers_0_probe_ready = ManagerTileLinkNetworkPort_2_io_manager_probe_ready;
  assign io_managers_0_release_valid = ManagerTileLinkNetworkPort_2_io_manager_release_valid;
  assign io_managers_0_release_bits_addr_beat = ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_beat;
  assign io_managers_0_release_bits_addr_block = ManagerTileLinkNetworkPort_2_io_manager_release_bits_addr_block;
  assign io_managers_0_release_bits_client_xact_id = ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_xact_id;
  assign io_managers_0_release_bits_voluntary = ManagerTileLinkNetworkPort_2_io_manager_release_bits_voluntary;
  assign io_managers_0_release_bits_r_type = ManagerTileLinkNetworkPort_2_io_manager_release_bits_r_type;
  assign io_managers_0_release_bits_data = ManagerTileLinkNetworkPort_2_io_manager_release_bits_data;
  assign io_managers_0_release_bits_client_id = ManagerTileLinkNetworkPort_2_io_manager_release_bits_client_id;
  assign io_managers_1_acquire_valid = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_valid;
  assign io_managers_1_acquire_bits_addr_block = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_block;
  assign io_managers_1_acquire_bits_client_xact_id = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_xact_id;
  assign io_managers_1_acquire_bits_addr_beat = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_addr_beat;
  assign io_managers_1_acquire_bits_is_builtin_type = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_is_builtin_type;
  assign io_managers_1_acquire_bits_a_type = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_a_type;
  assign io_managers_1_acquire_bits_union = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_union;
  assign io_managers_1_acquire_bits_data = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_data;
  assign io_managers_1_acquire_bits_client_id = ManagerTileLinkNetworkPort_1_1_io_manager_acquire_bits_client_id;
  assign io_managers_1_grant_ready = ManagerTileLinkNetworkPort_1_1_io_manager_grant_ready;
  assign io_managers_1_finish_valid = ManagerTileLinkNetworkPort_1_1_io_manager_finish_valid;
  assign io_managers_1_finish_bits_manager_xact_id = ManagerTileLinkNetworkPort_1_1_io_manager_finish_bits_manager_xact_id;
  assign io_managers_1_probe_ready = ManagerTileLinkNetworkPort_1_1_io_manager_probe_ready;
  assign io_managers_1_release_valid = ManagerTileLinkNetworkPort_1_1_io_manager_release_valid;
  assign io_managers_1_release_bits_addr_beat = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_beat;
  assign io_managers_1_release_bits_addr_block = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_addr_block;
  assign io_managers_1_release_bits_client_xact_id = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_xact_id;
  assign io_managers_1_release_bits_voluntary = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_voluntary;
  assign io_managers_1_release_bits_r_type = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_r_type;
  assign io_managers_1_release_bits_data = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_data;
  assign io_managers_1_release_bits_client_id = ManagerTileLinkNetworkPort_1_1_io_manager_release_bits_client_id;
  assign TileLinkEnqueuer_4_clk = clk;
  assign TileLinkEnqueuer_4_reset = reset;
  assign TileLinkEnqueuer_4_io_client_acquire_valid = ClientTileLinkNetworkPort_1_io_network_acquire_valid;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_header_src = ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_src;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_header_dst = ClientTileLinkNetworkPort_1_io_network_acquire_bits_header_dst;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_block = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_client_xact_id = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_addr_beat = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_is_builtin_type = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_a_type = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_union = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_union;
  assign TileLinkEnqueuer_4_io_client_acquire_bits_payload_data = ClientTileLinkNetworkPort_1_io_network_acquire_bits_payload_data;
  assign TileLinkEnqueuer_4_io_client_grant_ready = ClientTileLinkNetworkPort_1_io_network_grant_ready;
  assign TileLinkEnqueuer_4_io_client_finish_valid = ClientTileLinkNetworkPort_1_io_network_finish_valid;
  assign TileLinkEnqueuer_4_io_client_finish_bits_header_src = ClientTileLinkNetworkPort_1_io_network_finish_bits_header_src;
  assign TileLinkEnqueuer_4_io_client_finish_bits_header_dst = ClientTileLinkNetworkPort_1_io_network_finish_bits_header_dst;
  assign TileLinkEnqueuer_4_io_client_finish_bits_payload_manager_xact_id = ClientTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_4_io_client_probe_ready = ClientTileLinkNetworkPort_1_io_network_probe_ready;
  assign TileLinkEnqueuer_4_io_client_release_valid = ClientTileLinkNetworkPort_1_io_network_release_valid;
  assign TileLinkEnqueuer_4_io_client_release_bits_header_src = ClientTileLinkNetworkPort_1_io_network_release_bits_header_src;
  assign TileLinkEnqueuer_4_io_client_release_bits_header_dst = ClientTileLinkNetworkPort_1_io_network_release_bits_header_dst;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_addr_beat = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_addr_block = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_client_xact_id = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_voluntary = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_r_type = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_r_type;
  assign TileLinkEnqueuer_4_io_client_release_bits_payload_data = ClientTileLinkNetworkPort_1_io_network_release_bits_payload_data;
  assign TileLinkEnqueuer_4_io_manager_acquire_ready = T_13624_ready;
  assign TileLinkEnqueuer_4_io_manager_grant_valid = T_17371_valid;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_header_src = T_17371_bits_header_src;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_header_dst = T_17371_bits_header_dst;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_addr_beat = T_17371_bits_payload_addr_beat;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_client_xact_id = T_17371_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_manager_xact_id = T_17371_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_is_builtin_type = T_17371_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_g_type = T_17371_bits_payload_g_type;
  assign TileLinkEnqueuer_4_io_manager_grant_bits_payload_data = T_17371_bits_payload_data;
  assign TileLinkEnqueuer_4_io_manager_finish_ready = T_19326_ready;
  assign TileLinkEnqueuer_4_io_manager_probe_valid = T_15939_valid;
  assign TileLinkEnqueuer_4_io_manager_probe_bits_header_src = T_15939_bits_header_src;
  assign TileLinkEnqueuer_4_io_manager_probe_bits_header_dst = T_15939_bits_header_dst;
  assign TileLinkEnqueuer_4_io_manager_probe_bits_payload_addr_block = T_15939_bits_payload_addr_block;
  assign TileLinkEnqueuer_4_io_manager_probe_bits_payload_p_type = T_15939_bits_payload_p_type;
  assign TileLinkEnqueuer_4_io_manager_release_ready = T_15091_ready;
  assign ClientTileLinkNetworkPort_1_clk = clk;
  assign ClientTileLinkNetworkPort_1_reset = reset;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_valid = io_clients_cached_0_acquire_valid;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_block = io_clients_cached_0_acquire_bits_addr_block;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id = io_clients_cached_0_acquire_bits_client_xact_id;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat = io_clients_cached_0_acquire_bits_addr_beat;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type = io_clients_cached_0_acquire_bits_is_builtin_type;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_a_type = io_clients_cached_0_acquire_bits_a_type;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_union = io_clients_cached_0_acquire_bits_union;
  assign ClientTileLinkNetworkPort_1_io_client_acquire_bits_data = io_clients_cached_0_acquire_bits_data;
  assign ClientTileLinkNetworkPort_1_io_client_probe_ready = io_clients_cached_0_probe_ready;
  assign ClientTileLinkNetworkPort_1_io_client_release_valid = io_clients_cached_0_release_valid;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_addr_beat = io_clients_cached_0_release_bits_addr_beat;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_addr_block = io_clients_cached_0_release_bits_addr_block;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_client_xact_id = io_clients_cached_0_release_bits_client_xact_id;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_voluntary = io_clients_cached_0_release_bits_voluntary;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_r_type = io_clients_cached_0_release_bits_r_type;
  assign ClientTileLinkNetworkPort_1_io_client_release_bits_data = io_clients_cached_0_release_bits_data;
  assign ClientTileLinkNetworkPort_1_io_client_grant_ready = io_clients_cached_0_grant_ready;
  assign ClientTileLinkNetworkPort_1_io_client_finish_valid = io_clients_cached_0_finish_valid;
  assign ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_xact_id = io_clients_cached_0_finish_bits_manager_xact_id;
  assign ClientTileLinkNetworkPort_1_io_client_finish_bits_manager_id = io_clients_cached_0_finish_bits_manager_id;
  assign ClientTileLinkNetworkPort_1_io_network_acquire_ready = TileLinkEnqueuer_4_io_client_acquire_ready;
  assign ClientTileLinkNetworkPort_1_io_network_grant_valid = TileLinkEnqueuer_4_io_client_grant_valid;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_header_src = TileLinkEnqueuer_4_io_client_grant_bits_header_src;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_header_dst = TileLinkEnqueuer_4_io_client_grant_bits_header_dst;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat = TileLinkEnqueuer_4_io_client_grant_bits_payload_addr_beat;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id = TileLinkEnqueuer_4_io_client_grant_bits_payload_client_xact_id;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id = TileLinkEnqueuer_4_io_client_grant_bits_payload_manager_xact_id;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type = TileLinkEnqueuer_4_io_client_grant_bits_payload_is_builtin_type;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type = TileLinkEnqueuer_4_io_client_grant_bits_payload_g_type;
  assign ClientTileLinkNetworkPort_1_io_network_grant_bits_payload_data = TileLinkEnqueuer_4_io_client_grant_bits_payload_data;
  assign ClientTileLinkNetworkPort_1_io_network_finish_ready = TileLinkEnqueuer_4_io_client_finish_ready;
  assign ClientTileLinkNetworkPort_1_io_network_probe_valid = TileLinkEnqueuer_4_io_client_probe_valid;
  assign ClientTileLinkNetworkPort_1_io_network_probe_bits_header_src = TileLinkEnqueuer_4_io_client_probe_bits_header_src;
  assign ClientTileLinkNetworkPort_1_io_network_probe_bits_header_dst = TileLinkEnqueuer_4_io_client_probe_bits_header_dst;
  assign ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block = TileLinkEnqueuer_4_io_client_probe_bits_payload_addr_block;
  assign ClientTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type = TileLinkEnqueuer_4_io_client_probe_bits_payload_p_type;
  assign ClientTileLinkNetworkPort_1_io_network_release_ready = TileLinkEnqueuer_4_io_client_release_ready;
  assign TileLinkEnqueuer_1_1_clk = clk;
  assign TileLinkEnqueuer_1_1_reset = reset;
  assign TileLinkEnqueuer_1_1_io_client_acquire_valid = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_valid;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_header_src = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_src;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_header_dst = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_header_dst;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_block = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_block;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_client_xact_id = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_addr_beat = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_addr_beat;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_is_builtin_type = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_a_type = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_a_type;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_union = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_union;
  assign TileLinkEnqueuer_1_1_io_client_acquire_bits_payload_data = ClientUncachedTileLinkNetworkPort_1_io_network_acquire_bits_payload_data;
  assign TileLinkEnqueuer_1_1_io_client_grant_ready = ClientUncachedTileLinkNetworkPort_1_io_network_grant_ready;
  assign TileLinkEnqueuer_1_1_io_client_finish_valid = ClientUncachedTileLinkNetworkPort_1_io_network_finish_valid;
  assign TileLinkEnqueuer_1_1_io_client_finish_bits_header_src = ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_src;
  assign TileLinkEnqueuer_1_1_io_client_finish_bits_header_dst = ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_header_dst;
  assign TileLinkEnqueuer_1_1_io_client_finish_bits_payload_manager_xact_id = ClientUncachedTileLinkNetworkPort_1_io_network_finish_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_1_1_io_client_probe_ready = ClientUncachedTileLinkNetworkPort_1_io_network_probe_ready;
  assign TileLinkEnqueuer_1_1_io_client_release_valid = ClientUncachedTileLinkNetworkPort_1_io_network_release_valid;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_header_src = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_src;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_header_dst = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_header_dst;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_beat = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_beat;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_addr_block = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_addr_block;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_client_xact_id = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_voluntary = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_voluntary;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_r_type = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_r_type;
  assign TileLinkEnqueuer_1_1_io_client_release_bits_payload_data = ClientUncachedTileLinkNetworkPort_1_io_network_release_bits_payload_data;
  assign TileLinkEnqueuer_1_1_io_manager_acquire_ready = T_13794_ready;
  assign TileLinkEnqueuer_1_1_io_manager_grant_valid = T_17936_valid;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_header_src = T_17936_bits_header_src;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_header_dst = T_17936_bits_header_dst;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_addr_beat = T_17936_bits_payload_addr_beat;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_client_xact_id = T_17936_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_manager_xact_id = T_17936_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_is_builtin_type = T_17936_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_g_type = T_17936_bits_payload_g_type;
  assign TileLinkEnqueuer_1_1_io_manager_grant_bits_payload_data = T_17936_bits_payload_data;
  assign TileLinkEnqueuer_1_1_io_manager_finish_ready = T_19466_ready;
  assign TileLinkEnqueuer_1_1_io_manager_probe_valid = T_16484_valid;
  assign TileLinkEnqueuer_1_1_io_manager_probe_bits_header_src = T_16484_bits_header_src;
  assign TileLinkEnqueuer_1_1_io_manager_probe_bits_header_dst = T_16484_bits_header_dst;
  assign TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_addr_block = T_16484_bits_payload_addr_block;
  assign TileLinkEnqueuer_1_1_io_manager_probe_bits_payload_p_type = T_16484_bits_payload_p_type;
  assign TileLinkEnqueuer_1_1_io_manager_release_ready = T_15256_ready;
  assign ClientUncachedTileLinkNetworkPort_1_clk = clk;
  assign ClientUncachedTileLinkNetworkPort_1_reset = reset;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_valid = io_clients_uncached_0_acquire_valid;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_block = io_clients_uncached_0_acquire_bits_addr_block;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_client_xact_id = io_clients_uncached_0_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_addr_beat = io_clients_uncached_0_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_is_builtin_type = io_clients_uncached_0_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_a_type = io_clients_uncached_0_acquire_bits_a_type;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_union = io_clients_uncached_0_acquire_bits_union;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_acquire_bits_data = io_clients_uncached_0_acquire_bits_data;
  assign ClientUncachedTileLinkNetworkPort_1_io_client_grant_ready = io_clients_uncached_0_grant_ready;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_acquire_ready = TileLinkEnqueuer_1_1_io_client_acquire_ready;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_valid = TileLinkEnqueuer_1_1_io_client_grant_valid;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_src = TileLinkEnqueuer_1_1_io_client_grant_bits_header_src;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_header_dst = TileLinkEnqueuer_1_1_io_client_grant_bits_header_dst;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_addr_beat = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_addr_beat;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_client_xact_id = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_client_xact_id;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_manager_xact_id = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_manager_xact_id;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_is_builtin_type = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_is_builtin_type;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_g_type = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_g_type;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_grant_bits_payload_data = TileLinkEnqueuer_1_1_io_client_grant_bits_payload_data;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_finish_ready = TileLinkEnqueuer_1_1_io_client_finish_ready;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_probe_valid = TileLinkEnqueuer_1_1_io_client_probe_valid;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_src = TileLinkEnqueuer_1_1_io_client_probe_bits_header_src;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_header_dst = TileLinkEnqueuer_1_1_io_client_probe_bits_header_dst;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_addr_block = TileLinkEnqueuer_1_1_io_client_probe_bits_payload_addr_block;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_probe_bits_payload_p_type = TileLinkEnqueuer_1_1_io_client_probe_bits_payload_p_type;
  assign ClientUncachedTileLinkNetworkPort_1_io_network_release_ready = TileLinkEnqueuer_1_1_io_client_release_ready;
  assign ManagerTileLinkNetworkPort_2_clk = clk;
  assign ManagerTileLinkNetworkPort_2_reset = reset;
  assign ManagerTileLinkNetworkPort_2_io_manager_acquire_ready = io_managers_0_acquire_ready;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_valid = io_managers_0_grant_valid;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_addr_beat = io_managers_0_grant_bits_addr_beat;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_xact_id = io_managers_0_grant_bits_client_xact_id;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_manager_xact_id = io_managers_0_grant_bits_manager_xact_id;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_is_builtin_type = io_managers_0_grant_bits_is_builtin_type;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_g_type = io_managers_0_grant_bits_g_type;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_data = io_managers_0_grant_bits_data;
  assign ManagerTileLinkNetworkPort_2_io_manager_grant_bits_client_id = io_managers_0_grant_bits_client_id;
  assign ManagerTileLinkNetworkPort_2_io_manager_finish_ready = io_managers_0_finish_ready;
  assign ManagerTileLinkNetworkPort_2_io_manager_probe_valid = io_managers_0_probe_valid;
  assign ManagerTileLinkNetworkPort_2_io_manager_probe_bits_addr_block = io_managers_0_probe_bits_addr_block;
  assign ManagerTileLinkNetworkPort_2_io_manager_probe_bits_p_type = io_managers_0_probe_bits_p_type;
  assign ManagerTileLinkNetworkPort_2_io_manager_probe_bits_client_id = io_managers_0_probe_bits_client_id;
  assign ManagerTileLinkNetworkPort_2_io_manager_release_ready = io_managers_0_release_ready;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_valid = TileLinkEnqueuer_2_1_io_manager_acquire_valid;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_src = TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_src;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_header_dst = TileLinkEnqueuer_2_1_io_manager_acquire_bits_header_dst;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_block = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_block;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_client_xact_id = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_client_xact_id;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_addr_beat = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_addr_beat;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_is_builtin_type = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_is_builtin_type;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_a_type = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_a_type;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_union = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_union;
  assign ManagerTileLinkNetworkPort_2_io_network_acquire_bits_payload_data = TileLinkEnqueuer_2_1_io_manager_acquire_bits_payload_data;
  assign ManagerTileLinkNetworkPort_2_io_network_grant_ready = TileLinkEnqueuer_2_1_io_manager_grant_ready;
  assign ManagerTileLinkNetworkPort_2_io_network_finish_valid = TileLinkEnqueuer_2_1_io_manager_finish_valid;
  assign ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_src = TileLinkEnqueuer_2_1_io_manager_finish_bits_header_src;
  assign ManagerTileLinkNetworkPort_2_io_network_finish_bits_header_dst = TileLinkEnqueuer_2_1_io_manager_finish_bits_header_dst;
  assign ManagerTileLinkNetworkPort_2_io_network_finish_bits_payload_manager_xact_id = TileLinkEnqueuer_2_1_io_manager_finish_bits_payload_manager_xact_id;
  assign ManagerTileLinkNetworkPort_2_io_network_probe_ready = TileLinkEnqueuer_2_1_io_manager_probe_ready;
  assign ManagerTileLinkNetworkPort_2_io_network_release_valid = TileLinkEnqueuer_2_1_io_manager_release_valid;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_header_src = TileLinkEnqueuer_2_1_io_manager_release_bits_header_src;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_header_dst = TileLinkEnqueuer_2_1_io_manager_release_bits_header_dst;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_beat = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_beat;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_addr_block = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_addr_block;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_client_xact_id = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_client_xact_id;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_voluntary = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_voluntary;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_r_type = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_r_type;
  assign ManagerTileLinkNetworkPort_2_io_network_release_bits_payload_data = TileLinkEnqueuer_2_1_io_manager_release_bits_payload_data;
  assign TileLinkEnqueuer_2_1_clk = clk;
  assign TileLinkEnqueuer_2_1_reset = reset;
  assign TileLinkEnqueuer_2_1_io_client_acquire_valid = T_12724_valid;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_header_src = T_12724_bits_header_src;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_header_dst = T_12724_bits_header_dst;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_block = T_12724_bits_payload_addr_block;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_client_xact_id = T_12724_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_addr_beat = T_12724_bits_payload_addr_beat;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_is_builtin_type = T_12724_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_a_type = T_12724_bits_payload_a_type;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_union = T_12724_bits_payload_union;
  assign TileLinkEnqueuer_2_1_io_client_acquire_bits_payload_data = T_12724_bits_payload_data;
  assign TileLinkEnqueuer_2_1_io_client_grant_ready = T_16801_ready;
  assign TileLinkEnqueuer_2_1_io_client_finish_valid = T_18486_valid;
  assign TileLinkEnqueuer_2_1_io_client_finish_bits_header_src = T_18486_bits_header_src;
  assign TileLinkEnqueuer_2_1_io_client_finish_bits_header_dst = T_18486_bits_header_dst;
  assign TileLinkEnqueuer_2_1_io_client_finish_bits_payload_manager_xact_id = T_18486_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_2_1_io_client_probe_ready = T_15409_ready;
  assign TileLinkEnqueuer_2_1_io_client_release_valid = T_14201_valid;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_header_src = T_14201_bits_header_src;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_header_dst = T_14201_bits_header_dst;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_beat = T_14201_bits_payload_addr_beat;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_addr_block = T_14201_bits_payload_addr_block;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_client_xact_id = T_14201_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_voluntary = T_14201_bits_payload_voluntary;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_r_type = T_14201_bits_payload_r_type;
  assign TileLinkEnqueuer_2_1_io_client_release_bits_payload_data = T_14201_bits_payload_data;
  assign TileLinkEnqueuer_2_1_io_manager_acquire_ready = ManagerTileLinkNetworkPort_2_io_network_acquire_ready;
  assign TileLinkEnqueuer_2_1_io_manager_grant_valid = ManagerTileLinkNetworkPort_2_io_network_grant_valid;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_header_src = ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_src;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_header_dst = ManagerTileLinkNetworkPort_2_io_network_grant_bits_header_dst;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_addr_beat = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_addr_beat;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_client_xact_id = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_manager_xact_id = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_is_builtin_type = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_g_type = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_g_type;
  assign TileLinkEnqueuer_2_1_io_manager_grant_bits_payload_data = ManagerTileLinkNetworkPort_2_io_network_grant_bits_payload_data;
  assign TileLinkEnqueuer_2_1_io_manager_finish_ready = ManagerTileLinkNetworkPort_2_io_network_finish_ready;
  assign TileLinkEnqueuer_2_1_io_manager_probe_valid = ManagerTileLinkNetworkPort_2_io_network_probe_valid;
  assign TileLinkEnqueuer_2_1_io_manager_probe_bits_header_src = ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_src;
  assign TileLinkEnqueuer_2_1_io_manager_probe_bits_header_dst = ManagerTileLinkNetworkPort_2_io_network_probe_bits_header_dst;
  assign TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_addr_block = ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_addr_block;
  assign TileLinkEnqueuer_2_1_io_manager_probe_bits_payload_p_type = ManagerTileLinkNetworkPort_2_io_network_probe_bits_payload_p_type;
  assign TileLinkEnqueuer_2_1_io_manager_release_ready = ManagerTileLinkNetworkPort_2_io_network_release_ready;
  assign ManagerTileLinkNetworkPort_1_1_clk = clk;
  assign ManagerTileLinkNetworkPort_1_1_reset = reset;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_acquire_ready = io_managers_1_acquire_ready;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_valid = io_managers_1_grant_valid;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_addr_beat = io_managers_1_grant_bits_addr_beat;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_xact_id = io_managers_1_grant_bits_client_xact_id;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_manager_xact_id = io_managers_1_grant_bits_manager_xact_id;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_is_builtin_type = io_managers_1_grant_bits_is_builtin_type;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_g_type = io_managers_1_grant_bits_g_type;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_data = io_managers_1_grant_bits_data;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_grant_bits_client_id = io_managers_1_grant_bits_client_id;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_finish_ready = io_managers_1_finish_ready;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_probe_valid = io_managers_1_probe_valid;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_addr_block = io_managers_1_probe_bits_addr_block;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_p_type = io_managers_1_probe_bits_p_type;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_probe_bits_client_id = io_managers_1_probe_bits_client_id;
  assign ManagerTileLinkNetworkPort_1_1_io_manager_release_ready = io_managers_1_release_ready;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_valid = TileLinkEnqueuer_3_1_io_manager_acquire_valid;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_src = TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_src;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_header_dst = TileLinkEnqueuer_3_1_io_manager_acquire_bits_header_dst;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_block = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_block;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_client_xact_id = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_client_xact_id;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_addr_beat = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_addr_beat;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_is_builtin_type = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_is_builtin_type;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_a_type = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_a_type;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_union = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_union;
  assign ManagerTileLinkNetworkPort_1_1_io_network_acquire_bits_payload_data = TileLinkEnqueuer_3_1_io_manager_acquire_bits_payload_data;
  assign ManagerTileLinkNetworkPort_1_1_io_network_grant_ready = TileLinkEnqueuer_3_1_io_manager_grant_ready;
  assign ManagerTileLinkNetworkPort_1_1_io_network_finish_valid = TileLinkEnqueuer_3_1_io_manager_finish_valid;
  assign ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_src = TileLinkEnqueuer_3_1_io_manager_finish_bits_header_src;
  assign ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_header_dst = TileLinkEnqueuer_3_1_io_manager_finish_bits_header_dst;
  assign ManagerTileLinkNetworkPort_1_1_io_network_finish_bits_payload_manager_xact_id = TileLinkEnqueuer_3_1_io_manager_finish_bits_payload_manager_xact_id;
  assign ManagerTileLinkNetworkPort_1_1_io_network_probe_ready = TileLinkEnqueuer_3_1_io_manager_probe_ready;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_valid = TileLinkEnqueuer_3_1_io_manager_release_valid;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_src = TileLinkEnqueuer_3_1_io_manager_release_bits_header_src;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_header_dst = TileLinkEnqueuer_3_1_io_manager_release_bits_header_dst;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_beat = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_beat;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_addr_block = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_addr_block;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_client_xact_id = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_client_xact_id;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_voluntary = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_voluntary;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_r_type = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_r_type;
  assign ManagerTileLinkNetworkPort_1_1_io_network_release_bits_payload_data = TileLinkEnqueuer_3_1_io_manager_release_bits_payload_data;
  assign TileLinkEnqueuer_3_1_clk = clk;
  assign TileLinkEnqueuer_3_1_reset = reset;
  assign TileLinkEnqueuer_3_1_io_client_acquire_valid = T_13294_valid;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_header_src = T_13294_bits_header_src;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_header_dst = T_13294_bits_header_dst;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_block = T_13294_bits_payload_addr_block;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_client_xact_id = T_13294_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_addr_beat = T_13294_bits_payload_addr_beat;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_is_builtin_type = T_13294_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_a_type = T_13294_bits_payload_a_type;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_union = T_13294_bits_payload_union;
  assign TileLinkEnqueuer_3_1_io_client_acquire_bits_payload_data = T_13294_bits_payload_data;
  assign TileLinkEnqueuer_3_1_io_client_grant_ready = T_16966_ready;
  assign TileLinkEnqueuer_3_1_io_client_finish_valid = T_19026_valid;
  assign TileLinkEnqueuer_3_1_io_client_finish_bits_header_src = T_19026_bits_header_src;
  assign TileLinkEnqueuer_3_1_io_client_finish_bits_header_dst = T_19026_bits_header_dst;
  assign TileLinkEnqueuer_3_1_io_client_finish_bits_payload_manager_xact_id = T_19026_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_3_1_io_client_probe_ready = T_15554_ready;
  assign TileLinkEnqueuer_3_1_io_client_release_valid = T_14766_valid;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_header_src = T_14766_bits_header_src;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_header_dst = T_14766_bits_header_dst;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_beat = T_14766_bits_payload_addr_beat;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_addr_block = T_14766_bits_payload_addr_block;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_client_xact_id = T_14766_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_voluntary = T_14766_bits_payload_voluntary;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_r_type = T_14766_bits_payload_r_type;
  assign TileLinkEnqueuer_3_1_io_client_release_bits_payload_data = T_14766_bits_payload_data;
  assign TileLinkEnqueuer_3_1_io_manager_acquire_ready = ManagerTileLinkNetworkPort_1_1_io_network_acquire_ready;
  assign TileLinkEnqueuer_3_1_io_manager_grant_valid = ManagerTileLinkNetworkPort_1_1_io_network_grant_valid;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_header_src = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_src;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_header_dst = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_header_dst;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_addr_beat = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_addr_beat;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_client_xact_id = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_manager_xact_id = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_is_builtin_type = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_g_type = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_g_type;
  assign TileLinkEnqueuer_3_1_io_manager_grant_bits_payload_data = ManagerTileLinkNetworkPort_1_1_io_network_grant_bits_payload_data;
  assign TileLinkEnqueuer_3_1_io_manager_finish_ready = ManagerTileLinkNetworkPort_1_1_io_network_finish_ready;
  assign TileLinkEnqueuer_3_1_io_manager_probe_valid = ManagerTileLinkNetworkPort_1_1_io_network_probe_valid;
  assign TileLinkEnqueuer_3_1_io_manager_probe_bits_header_src = ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_src;
  assign TileLinkEnqueuer_3_1_io_manager_probe_bits_header_dst = ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_header_dst;
  assign TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_addr_block = ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_addr_block;
  assign TileLinkEnqueuer_3_1_io_manager_probe_bits_payload_p_type = ManagerTileLinkNetworkPort_1_1_io_network_probe_bits_payload_p_type;
  assign TileLinkEnqueuer_3_1_io_manager_release_ready = ManagerTileLinkNetworkPort_1_1_io_network_release_ready;
  assign acqNet_clk = clk;
  assign acqNet_reset = reset;
  assign acqNet_io_in_0_valid = 1'h0;
  assign acqNet_io_in_0_bits_header_src = GEN_0;
  assign acqNet_io_in_0_bits_header_dst = GEN_1;
  assign acqNet_io_in_0_bits_payload_addr_block = GEN_2;
  assign acqNet_io_in_0_bits_payload_client_xact_id = GEN_3;
  assign acqNet_io_in_0_bits_payload_addr_beat = GEN_4;
  assign acqNet_io_in_0_bits_payload_is_builtin_type = GEN_5;
  assign acqNet_io_in_0_bits_payload_a_type = GEN_6;
  assign acqNet_io_in_0_bits_payload_union = GEN_7;
  assign acqNet_io_in_0_bits_payload_data = GEN_8;
  assign acqNet_io_in_1_valid = 1'h0;
  assign acqNet_io_in_1_bits_header_src = GEN_9;
  assign acqNet_io_in_1_bits_header_dst = GEN_10;
  assign acqNet_io_in_1_bits_payload_addr_block = GEN_11;
  assign acqNet_io_in_1_bits_payload_client_xact_id = GEN_12;
  assign acqNet_io_in_1_bits_payload_addr_beat = GEN_13;
  assign acqNet_io_in_1_bits_payload_is_builtin_type = GEN_14;
  assign acqNet_io_in_1_bits_payload_a_type = GEN_15;
  assign acqNet_io_in_1_bits_payload_union = GEN_16;
  assign acqNet_io_in_1_bits_payload_data = GEN_17;
  assign acqNet_io_in_2_valid = T_13624_valid;
  assign acqNet_io_in_2_bits_header_src = T_13624_bits_header_src;
  assign acqNet_io_in_2_bits_header_dst = T_13624_bits_header_dst;
  assign acqNet_io_in_2_bits_payload_addr_block = T_13624_bits_payload_addr_block;
  assign acqNet_io_in_2_bits_payload_client_xact_id = T_13624_bits_payload_client_xact_id;
  assign acqNet_io_in_2_bits_payload_addr_beat = T_13624_bits_payload_addr_beat;
  assign acqNet_io_in_2_bits_payload_is_builtin_type = T_13624_bits_payload_is_builtin_type;
  assign acqNet_io_in_2_bits_payload_a_type = T_13624_bits_payload_a_type;
  assign acqNet_io_in_2_bits_payload_union = T_13624_bits_payload_union;
  assign acqNet_io_in_2_bits_payload_data = T_13624_bits_payload_data;
  assign acqNet_io_in_3_valid = T_13794_valid;
  assign acqNet_io_in_3_bits_header_src = T_13794_bits_header_src;
  assign acqNet_io_in_3_bits_header_dst = T_13794_bits_header_dst;
  assign acqNet_io_in_3_bits_payload_addr_block = T_13794_bits_payload_addr_block;
  assign acqNet_io_in_3_bits_payload_client_xact_id = T_13794_bits_payload_client_xact_id;
  assign acqNet_io_in_3_bits_payload_addr_beat = T_13794_bits_payload_addr_beat;
  assign acqNet_io_in_3_bits_payload_is_builtin_type = T_13794_bits_payload_is_builtin_type;
  assign acqNet_io_in_3_bits_payload_a_type = T_13794_bits_payload_a_type;
  assign acqNet_io_in_3_bits_payload_union = T_13794_bits_payload_union;
  assign acqNet_io_in_3_bits_payload_data = T_13794_bits_payload_data;
  assign acqNet_io_out_0_ready = T_12724_ready;
  assign acqNet_io_out_1_ready = T_13294_ready;
  assign acqNet_io_out_2_ready = 1'h0;
  assign acqNet_io_out_3_ready = 1'h0;
  assign relNet_clk = clk;
  assign relNet_reset = reset;
  assign relNet_io_in_0_valid = 1'h0;
  assign relNet_io_in_0_bits_header_src = GEN_18;
  assign relNet_io_in_0_bits_header_dst = GEN_19;
  assign relNet_io_in_0_bits_payload_addr_beat = GEN_20;
  assign relNet_io_in_0_bits_payload_addr_block = GEN_21;
  assign relNet_io_in_0_bits_payload_client_xact_id = GEN_22;
  assign relNet_io_in_0_bits_payload_voluntary = GEN_23;
  assign relNet_io_in_0_bits_payload_r_type = GEN_24;
  assign relNet_io_in_0_bits_payload_data = GEN_25;
  assign relNet_io_in_1_valid = 1'h0;
  assign relNet_io_in_1_bits_header_src = GEN_26;
  assign relNet_io_in_1_bits_header_dst = GEN_27;
  assign relNet_io_in_1_bits_payload_addr_beat = GEN_28;
  assign relNet_io_in_1_bits_payload_addr_block = GEN_29;
  assign relNet_io_in_1_bits_payload_client_xact_id = GEN_30;
  assign relNet_io_in_1_bits_payload_voluntary = GEN_31;
  assign relNet_io_in_1_bits_payload_r_type = GEN_32;
  assign relNet_io_in_1_bits_payload_data = GEN_33;
  assign relNet_io_in_2_valid = T_15091_valid;
  assign relNet_io_in_2_bits_header_src = T_15091_bits_header_src;
  assign relNet_io_in_2_bits_header_dst = T_15091_bits_header_dst;
  assign relNet_io_in_2_bits_payload_addr_beat = T_15091_bits_payload_addr_beat;
  assign relNet_io_in_2_bits_payload_addr_block = T_15091_bits_payload_addr_block;
  assign relNet_io_in_2_bits_payload_client_xact_id = T_15091_bits_payload_client_xact_id;
  assign relNet_io_in_2_bits_payload_voluntary = T_15091_bits_payload_voluntary;
  assign relNet_io_in_2_bits_payload_r_type = T_15091_bits_payload_r_type;
  assign relNet_io_in_2_bits_payload_data = T_15091_bits_payload_data;
  assign relNet_io_in_3_valid = T_15256_valid;
  assign relNet_io_in_3_bits_header_src = T_15256_bits_header_src;
  assign relNet_io_in_3_bits_header_dst = T_15256_bits_header_dst;
  assign relNet_io_in_3_bits_payload_addr_beat = T_15256_bits_payload_addr_beat;
  assign relNet_io_in_3_bits_payload_addr_block = T_15256_bits_payload_addr_block;
  assign relNet_io_in_3_bits_payload_client_xact_id = T_15256_bits_payload_client_xact_id;
  assign relNet_io_in_3_bits_payload_voluntary = T_15256_bits_payload_voluntary;
  assign relNet_io_in_3_bits_payload_r_type = T_15256_bits_payload_r_type;
  assign relNet_io_in_3_bits_payload_data = T_15256_bits_payload_data;
  assign relNet_io_out_0_ready = T_14201_ready;
  assign relNet_io_out_1_ready = T_14766_ready;
  assign relNet_io_out_2_ready = 1'h0;
  assign relNet_io_out_3_ready = 1'h0;
  assign prbNet_clk = clk;
  assign prbNet_reset = reset;
  assign prbNet_io_in_0_valid = T_15409_valid;
  assign prbNet_io_in_0_bits_header_src = T_15409_bits_header_src;
  assign prbNet_io_in_0_bits_header_dst = T_15409_bits_header_dst;
  assign prbNet_io_in_0_bits_payload_addr_block = T_15409_bits_payload_addr_block;
  assign prbNet_io_in_0_bits_payload_p_type = T_15409_bits_payload_p_type;
  assign prbNet_io_in_1_valid = T_15554_valid;
  assign prbNet_io_in_1_bits_header_src = T_15554_bits_header_src;
  assign prbNet_io_in_1_bits_header_dst = T_15554_bits_header_dst;
  assign prbNet_io_in_1_bits_payload_addr_block = T_15554_bits_payload_addr_block;
  assign prbNet_io_in_1_bits_payload_p_type = T_15554_bits_payload_p_type;
  assign prbNet_io_in_2_valid = 1'h0;
  assign prbNet_io_in_2_bits_header_src = GEN_34;
  assign prbNet_io_in_2_bits_header_dst = GEN_35;
  assign prbNet_io_in_2_bits_payload_addr_block = GEN_36;
  assign prbNet_io_in_2_bits_payload_p_type = GEN_37;
  assign prbNet_io_in_3_valid = 1'h0;
  assign prbNet_io_in_3_bits_header_src = GEN_38;
  assign prbNet_io_in_3_bits_header_dst = GEN_39;
  assign prbNet_io_in_3_bits_payload_addr_block = GEN_40;
  assign prbNet_io_in_3_bits_payload_p_type = GEN_41;
  assign prbNet_io_out_0_ready = 1'h0;
  assign prbNet_io_out_1_ready = 1'h0;
  assign prbNet_io_out_2_ready = T_15939_ready;
  assign prbNet_io_out_3_ready = T_16484_ready;
  assign gntNet_clk = clk;
  assign gntNet_reset = reset;
  assign gntNet_io_in_0_valid = T_16801_valid;
  assign gntNet_io_in_0_bits_header_src = T_16801_bits_header_src;
  assign gntNet_io_in_0_bits_header_dst = T_16801_bits_header_dst;
  assign gntNet_io_in_0_bits_payload_addr_beat = T_16801_bits_payload_addr_beat;
  assign gntNet_io_in_0_bits_payload_client_xact_id = T_16801_bits_payload_client_xact_id;
  assign gntNet_io_in_0_bits_payload_manager_xact_id = T_16801_bits_payload_manager_xact_id;
  assign gntNet_io_in_0_bits_payload_is_builtin_type = T_16801_bits_payload_is_builtin_type;
  assign gntNet_io_in_0_bits_payload_g_type = T_16801_bits_payload_g_type;
  assign gntNet_io_in_0_bits_payload_data = T_16801_bits_payload_data;
  assign gntNet_io_in_1_valid = T_16966_valid;
  assign gntNet_io_in_1_bits_header_src = T_16966_bits_header_src;
  assign gntNet_io_in_1_bits_header_dst = T_16966_bits_header_dst;
  assign gntNet_io_in_1_bits_payload_addr_beat = T_16966_bits_payload_addr_beat;
  assign gntNet_io_in_1_bits_payload_client_xact_id = T_16966_bits_payload_client_xact_id;
  assign gntNet_io_in_1_bits_payload_manager_xact_id = T_16966_bits_payload_manager_xact_id;
  assign gntNet_io_in_1_bits_payload_is_builtin_type = T_16966_bits_payload_is_builtin_type;
  assign gntNet_io_in_1_bits_payload_g_type = T_16966_bits_payload_g_type;
  assign gntNet_io_in_1_bits_payload_data = T_16966_bits_payload_data;
  assign gntNet_io_in_2_valid = 1'h0;
  assign gntNet_io_in_2_bits_header_src = GEN_42;
  assign gntNet_io_in_2_bits_header_dst = GEN_43;
  assign gntNet_io_in_2_bits_payload_addr_beat = GEN_44;
  assign gntNet_io_in_2_bits_payload_client_xact_id = GEN_45;
  assign gntNet_io_in_2_bits_payload_manager_xact_id = GEN_46;
  assign gntNet_io_in_2_bits_payload_is_builtin_type = GEN_47;
  assign gntNet_io_in_2_bits_payload_g_type = GEN_48;
  assign gntNet_io_in_2_bits_payload_data = GEN_49;
  assign gntNet_io_in_3_valid = 1'h0;
  assign gntNet_io_in_3_bits_header_src = GEN_50;
  assign gntNet_io_in_3_bits_header_dst = GEN_51;
  assign gntNet_io_in_3_bits_payload_addr_beat = GEN_52;
  assign gntNet_io_in_3_bits_payload_client_xact_id = GEN_53;
  assign gntNet_io_in_3_bits_payload_manager_xact_id = GEN_54;
  assign gntNet_io_in_3_bits_payload_is_builtin_type = GEN_55;
  assign gntNet_io_in_3_bits_payload_g_type = GEN_56;
  assign gntNet_io_in_3_bits_payload_data = GEN_57;
  assign gntNet_io_out_0_ready = 1'h0;
  assign gntNet_io_out_1_ready = 1'h0;
  assign gntNet_io_out_2_ready = T_17371_ready;
  assign gntNet_io_out_3_ready = T_17936_ready;
  assign ackNet_clk = clk;
  assign ackNet_reset = reset;
  assign ackNet_io_in_0_valid = 1'h0;
  assign ackNet_io_in_0_bits_header_src = GEN_58;
  assign ackNet_io_in_0_bits_header_dst = GEN_59;
  assign ackNet_io_in_0_bits_payload_manager_xact_id = GEN_60;
  assign ackNet_io_in_1_valid = 1'h0;
  assign ackNet_io_in_1_bits_header_src = GEN_61;
  assign ackNet_io_in_1_bits_header_dst = GEN_62;
  assign ackNet_io_in_1_bits_payload_manager_xact_id = GEN_63;
  assign ackNet_io_in_2_valid = T_19326_valid;
  assign ackNet_io_in_2_bits_header_src = T_19326_bits_header_src;
  assign ackNet_io_in_2_bits_header_dst = T_19326_bits_header_dst;
  assign ackNet_io_in_2_bits_payload_manager_xact_id = T_19326_bits_payload_manager_xact_id;
  assign ackNet_io_in_3_valid = T_19466_valid;
  assign ackNet_io_in_3_bits_header_src = T_19466_bits_header_src;
  assign ackNet_io_in_3_bits_header_dst = T_19466_bits_header_dst;
  assign ackNet_io_in_3_bits_payload_manager_xact_id = T_19466_bits_payload_manager_xact_id;
  assign ackNet_io_out_0_ready = T_18486_ready;
  assign ackNet_io_out_1_ready = T_19026_ready;
  assign ackNet_io_out_2_ready = 1'h0;
  assign ackNet_io_out_3_ready = 1'h0;
  assign T_12724_ready = TileLinkEnqueuer_2_1_io_client_acquire_ready;
  assign T_12724_valid = acqNet_io_out_0_valid;
  assign T_12724_bits_header_src = T_12953;
  assign T_12724_bits_header_dst = acqNet_io_out_0_bits_header_dst;
  assign T_12724_bits_payload_addr_block = acqNet_io_out_0_bits_payload_addr_block;
  assign T_12724_bits_payload_client_xact_id = acqNet_io_out_0_bits_payload_client_xact_id;
  assign T_12724_bits_payload_addr_beat = acqNet_io_out_0_bits_payload_addr_beat;
  assign T_12724_bits_payload_is_builtin_type = acqNet_io_out_0_bits_payload_is_builtin_type;
  assign T_12724_bits_payload_a_type = acqNet_io_out_0_bits_payload_a_type;
  assign T_12724_bits_payload_union = acqNet_io_out_0_bits_payload_union;
  assign T_12724_bits_payload_data = acqNet_io_out_0_bits_payload_data;
  assign T_12952 = acqNet_io_out_0_bits_header_src - 2'h2;
  assign T_12953 = T_12952[1:0];
  assign T_13294_ready = TileLinkEnqueuer_3_1_io_client_acquire_ready;
  assign T_13294_valid = acqNet_io_out_1_valid;
  assign T_13294_bits_header_src = T_13523;
  assign T_13294_bits_header_dst = acqNet_io_out_1_bits_header_dst;
  assign T_13294_bits_payload_addr_block = acqNet_io_out_1_bits_payload_addr_block;
  assign T_13294_bits_payload_client_xact_id = acqNet_io_out_1_bits_payload_client_xact_id;
  assign T_13294_bits_payload_addr_beat = acqNet_io_out_1_bits_payload_addr_beat;
  assign T_13294_bits_payload_is_builtin_type = acqNet_io_out_1_bits_payload_is_builtin_type;
  assign T_13294_bits_payload_a_type = acqNet_io_out_1_bits_payload_a_type;
  assign T_13294_bits_payload_union = acqNet_io_out_1_bits_payload_union;
  assign T_13294_bits_payload_data = acqNet_io_out_1_bits_payload_data;
  assign T_13522 = acqNet_io_out_1_bits_header_src - 2'h2;
  assign T_13523 = T_13522[1:0];
  assign T_13624_ready = acqNet_io_in_2_ready;
  assign T_13624_valid = TileLinkEnqueuer_4_io_manager_acquire_valid;
  assign T_13624_bits_header_src = T_13693;
  assign T_13624_bits_header_dst = TileLinkEnqueuer_4_io_manager_acquire_bits_header_dst;
  assign T_13624_bits_payload_addr_block = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_block;
  assign T_13624_bits_payload_client_xact_id = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_client_xact_id;
  assign T_13624_bits_payload_addr_beat = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_addr_beat;
  assign T_13624_bits_payload_is_builtin_type = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_is_builtin_type;
  assign T_13624_bits_payload_a_type = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_a_type;
  assign T_13624_bits_payload_union = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_union;
  assign T_13624_bits_payload_data = TileLinkEnqueuer_4_io_manager_acquire_bits_payload_data;
  assign T_13692 = TileLinkEnqueuer_4_io_manager_acquire_bits_header_src + 2'h2;
  assign T_13693 = T_13692[1:0];
  assign T_13794_ready = acqNet_io_in_3_ready;
  assign T_13794_valid = TileLinkEnqueuer_1_1_io_manager_acquire_valid;
  assign T_13794_bits_header_src = T_13863;
  assign T_13794_bits_header_dst = TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_dst;
  assign T_13794_bits_payload_addr_block = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_block;
  assign T_13794_bits_payload_client_xact_id = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_client_xact_id;
  assign T_13794_bits_payload_addr_beat = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_addr_beat;
  assign T_13794_bits_payload_is_builtin_type = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_is_builtin_type;
  assign T_13794_bits_payload_a_type = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_a_type;
  assign T_13794_bits_payload_union = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_union;
  assign T_13794_bits_payload_data = TileLinkEnqueuer_1_1_io_manager_acquire_bits_payload_data;
  assign T_13862 = TileLinkEnqueuer_1_1_io_manager_acquire_bits_header_src + 2'h2;
  assign T_13863 = T_13862[1:0];
  assign T_14201_ready = TileLinkEnqueuer_2_1_io_client_release_ready;
  assign T_14201_valid = relNet_io_out_0_valid;
  assign T_14201_bits_header_src = T_14428;
  assign T_14201_bits_header_dst = relNet_io_out_0_bits_header_dst;
  assign T_14201_bits_payload_addr_beat = relNet_io_out_0_bits_payload_addr_beat;
  assign T_14201_bits_payload_addr_block = relNet_io_out_0_bits_payload_addr_block;
  assign T_14201_bits_payload_client_xact_id = relNet_io_out_0_bits_payload_client_xact_id;
  assign T_14201_bits_payload_voluntary = relNet_io_out_0_bits_payload_voluntary;
  assign T_14201_bits_payload_r_type = relNet_io_out_0_bits_payload_r_type;
  assign T_14201_bits_payload_data = relNet_io_out_0_bits_payload_data;
  assign T_14427 = relNet_io_out_0_bits_header_src - 2'h2;
  assign T_14428 = T_14427[1:0];
  assign T_14766_ready = TileLinkEnqueuer_3_1_io_client_release_ready;
  assign T_14766_valid = relNet_io_out_1_valid;
  assign T_14766_bits_header_src = T_14993;
  assign T_14766_bits_header_dst = relNet_io_out_1_bits_header_dst;
  assign T_14766_bits_payload_addr_beat = relNet_io_out_1_bits_payload_addr_beat;
  assign T_14766_bits_payload_addr_block = relNet_io_out_1_bits_payload_addr_block;
  assign T_14766_bits_payload_client_xact_id = relNet_io_out_1_bits_payload_client_xact_id;
  assign T_14766_bits_payload_voluntary = relNet_io_out_1_bits_payload_voluntary;
  assign T_14766_bits_payload_r_type = relNet_io_out_1_bits_payload_r_type;
  assign T_14766_bits_payload_data = relNet_io_out_1_bits_payload_data;
  assign T_14992 = relNet_io_out_1_bits_header_src - 2'h2;
  assign T_14993 = T_14992[1:0];
  assign T_15091_ready = relNet_io_in_2_ready;
  assign T_15091_valid = TileLinkEnqueuer_4_io_manager_release_valid;
  assign T_15091_bits_header_src = T_15158;
  assign T_15091_bits_header_dst = TileLinkEnqueuer_4_io_manager_release_bits_header_dst;
  assign T_15091_bits_payload_addr_beat = TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_beat;
  assign T_15091_bits_payload_addr_block = TileLinkEnqueuer_4_io_manager_release_bits_payload_addr_block;
  assign T_15091_bits_payload_client_xact_id = TileLinkEnqueuer_4_io_manager_release_bits_payload_client_xact_id;
  assign T_15091_bits_payload_voluntary = TileLinkEnqueuer_4_io_manager_release_bits_payload_voluntary;
  assign T_15091_bits_payload_r_type = TileLinkEnqueuer_4_io_manager_release_bits_payload_r_type;
  assign T_15091_bits_payload_data = TileLinkEnqueuer_4_io_manager_release_bits_payload_data;
  assign T_15157 = TileLinkEnqueuer_4_io_manager_release_bits_header_src + 2'h2;
  assign T_15158 = T_15157[1:0];
  assign T_15256_ready = relNet_io_in_3_ready;
  assign T_15256_valid = TileLinkEnqueuer_1_1_io_manager_release_valid;
  assign T_15256_bits_header_src = T_15323;
  assign T_15256_bits_header_dst = TileLinkEnqueuer_1_1_io_manager_release_bits_header_dst;
  assign T_15256_bits_payload_addr_beat = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_beat;
  assign T_15256_bits_payload_addr_block = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_addr_block;
  assign T_15256_bits_payload_client_xact_id = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_client_xact_id;
  assign T_15256_bits_payload_voluntary = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_voluntary;
  assign T_15256_bits_payload_r_type = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_r_type;
  assign T_15256_bits_payload_data = TileLinkEnqueuer_1_1_io_manager_release_bits_payload_data;
  assign T_15322 = TileLinkEnqueuer_1_1_io_manager_release_bits_header_src + 2'h2;
  assign T_15323 = T_15322[1:0];
  assign T_15409_ready = prbNet_io_in_0_ready;
  assign T_15409_valid = TileLinkEnqueuer_2_1_io_client_probe_valid;
  assign T_15409_bits_header_src = TileLinkEnqueuer_2_1_io_client_probe_bits_header_src;
  assign T_15409_bits_header_dst = T_15468;
  assign T_15409_bits_payload_addr_block = TileLinkEnqueuer_2_1_io_client_probe_bits_payload_addr_block;
  assign T_15409_bits_payload_p_type = TileLinkEnqueuer_2_1_io_client_probe_bits_payload_p_type;
  assign T_15467 = TileLinkEnqueuer_2_1_io_client_probe_bits_header_dst + 2'h2;
  assign T_15468 = T_15467[1:0];
  assign T_15554_ready = prbNet_io_in_1_ready;
  assign T_15554_valid = TileLinkEnqueuer_3_1_io_client_probe_valid;
  assign T_15554_bits_header_src = TileLinkEnqueuer_3_1_io_client_probe_bits_header_src;
  assign T_15554_bits_header_dst = T_15613;
  assign T_15554_bits_payload_addr_block = TileLinkEnqueuer_3_1_io_client_probe_bits_payload_addr_block;
  assign T_15554_bits_payload_p_type = TileLinkEnqueuer_3_1_io_client_probe_bits_payload_p_type;
  assign T_15612 = TileLinkEnqueuer_3_1_io_client_probe_bits_header_dst + 2'h2;
  assign T_15613 = T_15612[1:0];
  assign T_15939_ready = TileLinkEnqueuer_4_io_manager_probe_ready;
  assign T_15939_valid = prbNet_io_out_2_valid;
  assign T_15939_bits_header_src = prbNet_io_out_2_bits_header_src;
  assign T_15939_bits_header_dst = T_16158;
  assign T_15939_bits_payload_addr_block = prbNet_io_out_2_bits_payload_addr_block;
  assign T_15939_bits_payload_p_type = prbNet_io_out_2_bits_payload_p_type;
  assign T_16157 = prbNet_io_out_2_bits_header_dst - 2'h2;
  assign T_16158 = T_16157[1:0];
  assign T_16484_ready = TileLinkEnqueuer_1_1_io_manager_probe_ready;
  assign T_16484_valid = prbNet_io_out_3_valid;
  assign T_16484_bits_header_src = prbNet_io_out_3_bits_header_src;
  assign T_16484_bits_header_dst = T_16703;
  assign T_16484_bits_payload_addr_block = prbNet_io_out_3_bits_payload_addr_block;
  assign T_16484_bits_payload_p_type = prbNet_io_out_3_bits_payload_p_type;
  assign T_16702 = prbNet_io_out_3_bits_header_dst - 2'h2;
  assign T_16703 = T_16702[1:0];
  assign T_16801_ready = gntNet_io_in_0_ready;
  assign T_16801_valid = TileLinkEnqueuer_2_1_io_client_grant_valid;
  assign T_16801_bits_header_src = TileLinkEnqueuer_2_1_io_client_grant_bits_header_src;
  assign T_16801_bits_header_dst = T_16868;
  assign T_16801_bits_payload_addr_beat = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_addr_beat;
  assign T_16801_bits_payload_client_xact_id = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_client_xact_id;
  assign T_16801_bits_payload_manager_xact_id = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_manager_xact_id;
  assign T_16801_bits_payload_is_builtin_type = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_is_builtin_type;
  assign T_16801_bits_payload_g_type = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_g_type;
  assign T_16801_bits_payload_data = TileLinkEnqueuer_2_1_io_client_grant_bits_payload_data;
  assign T_16867 = TileLinkEnqueuer_2_1_io_client_grant_bits_header_dst + 2'h2;
  assign T_16868 = T_16867[1:0];
  assign T_16966_ready = gntNet_io_in_1_ready;
  assign T_16966_valid = TileLinkEnqueuer_3_1_io_client_grant_valid;
  assign T_16966_bits_header_src = TileLinkEnqueuer_3_1_io_client_grant_bits_header_src;
  assign T_16966_bits_header_dst = T_17033;
  assign T_16966_bits_payload_addr_beat = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_addr_beat;
  assign T_16966_bits_payload_client_xact_id = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_client_xact_id;
  assign T_16966_bits_payload_manager_xact_id = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_manager_xact_id;
  assign T_16966_bits_payload_is_builtin_type = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_is_builtin_type;
  assign T_16966_bits_payload_g_type = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_g_type;
  assign T_16966_bits_payload_data = TileLinkEnqueuer_3_1_io_client_grant_bits_payload_data;
  assign T_17032 = TileLinkEnqueuer_3_1_io_client_grant_bits_header_dst + 2'h2;
  assign T_17033 = T_17032[1:0];
  assign T_17371_ready = TileLinkEnqueuer_4_io_manager_grant_ready;
  assign T_17371_valid = gntNet_io_out_2_valid;
  assign T_17371_bits_header_src = gntNet_io_out_2_bits_header_src;
  assign T_17371_bits_header_dst = T_17598;
  assign T_17371_bits_payload_addr_beat = gntNet_io_out_2_bits_payload_addr_beat;
  assign T_17371_bits_payload_client_xact_id = gntNet_io_out_2_bits_payload_client_xact_id;
  assign T_17371_bits_payload_manager_xact_id = gntNet_io_out_2_bits_payload_manager_xact_id;
  assign T_17371_bits_payload_is_builtin_type = gntNet_io_out_2_bits_payload_is_builtin_type;
  assign T_17371_bits_payload_g_type = gntNet_io_out_2_bits_payload_g_type;
  assign T_17371_bits_payload_data = gntNet_io_out_2_bits_payload_data;
  assign T_17597 = gntNet_io_out_2_bits_header_dst - 2'h2;
  assign T_17598 = T_17597[1:0];
  assign T_17936_ready = TileLinkEnqueuer_1_1_io_manager_grant_ready;
  assign T_17936_valid = gntNet_io_out_3_valid;
  assign T_17936_bits_header_src = gntNet_io_out_3_bits_header_src;
  assign T_17936_bits_header_dst = T_18163;
  assign T_17936_bits_payload_addr_beat = gntNet_io_out_3_bits_payload_addr_beat;
  assign T_17936_bits_payload_client_xact_id = gntNet_io_out_3_bits_payload_client_xact_id;
  assign T_17936_bits_payload_manager_xact_id = gntNet_io_out_3_bits_payload_manager_xact_id;
  assign T_17936_bits_payload_is_builtin_type = gntNet_io_out_3_bits_payload_is_builtin_type;
  assign T_17936_bits_payload_g_type = gntNet_io_out_3_bits_payload_g_type;
  assign T_17936_bits_payload_data = gntNet_io_out_3_bits_payload_data;
  assign T_18162 = gntNet_io_out_3_bits_header_dst - 2'h2;
  assign T_18163 = T_18162[1:0];
  assign T_18486_ready = TileLinkEnqueuer_2_1_io_client_finish_ready;
  assign T_18486_valid = ackNet_io_out_0_valid;
  assign T_18486_bits_header_src = T_18703;
  assign T_18486_bits_header_dst = ackNet_io_out_0_bits_header_dst;
  assign T_18486_bits_payload_manager_xact_id = ackNet_io_out_0_bits_payload_manager_xact_id;
  assign T_18702 = ackNet_io_out_0_bits_header_src - 2'h2;
  assign T_18703 = T_18702[1:0];
  assign T_19026_ready = TileLinkEnqueuer_3_1_io_client_finish_ready;
  assign T_19026_valid = ackNet_io_out_1_valid;
  assign T_19026_bits_header_src = T_19243;
  assign T_19026_bits_header_dst = ackNet_io_out_1_bits_header_dst;
  assign T_19026_bits_payload_manager_xact_id = ackNet_io_out_1_bits_payload_manager_xact_id;
  assign T_19242 = ackNet_io_out_1_bits_header_src - 2'h2;
  assign T_19243 = T_19242[1:0];
  assign T_19326_ready = ackNet_io_in_2_ready;
  assign T_19326_valid = TileLinkEnqueuer_4_io_manager_finish_valid;
  assign T_19326_bits_header_src = T_19383;
  assign T_19326_bits_header_dst = TileLinkEnqueuer_4_io_manager_finish_bits_header_dst;
  assign T_19326_bits_payload_manager_xact_id = TileLinkEnqueuer_4_io_manager_finish_bits_payload_manager_xact_id;
  assign T_19382 = TileLinkEnqueuer_4_io_manager_finish_bits_header_src + 2'h2;
  assign T_19383 = T_19382[1:0];
  assign T_19466_ready = ackNet_io_in_3_ready;
  assign T_19466_valid = TileLinkEnqueuer_1_1_io_manager_finish_valid;
  assign T_19466_bits_header_src = T_19523;
  assign T_19466_bits_header_dst = TileLinkEnqueuer_1_1_io_manager_finish_bits_header_dst;
  assign T_19466_bits_payload_manager_xact_id = TileLinkEnqueuer_1_1_io_manager_finish_bits_payload_manager_xact_id;
  assign T_19522 = TileLinkEnqueuer_1_1_io_manager_finish_bits_header_src + 2'h2;
  assign T_19523 = T_19522[1:0];
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_64 = {1{$random}};
  GEN_0 = GEN_64[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_65 = {1{$random}};
  GEN_1 = GEN_65[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_66 = {1{$random}};
  GEN_2 = GEN_66[25:0];
  `endif
  `ifdef RANDOMIZE
  GEN_67 = {1{$random}};
  GEN_3 = GEN_67[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_68 = {1{$random}};
  GEN_4 = GEN_68[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_69 = {1{$random}};
  GEN_5 = GEN_69[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_70 = {1{$random}};
  GEN_6 = GEN_70[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_71 = {1{$random}};
  GEN_7 = GEN_71[11:0];
  `endif
  `ifdef RANDOMIZE
  GEN_72 = {2{$random}};
  GEN_8 = GEN_72[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_73 = {1{$random}};
  GEN_9 = GEN_73[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_74 = {1{$random}};
  GEN_10 = GEN_74[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_75 = {1{$random}};
  GEN_11 = GEN_75[25:0];
  `endif
  `ifdef RANDOMIZE
  GEN_76 = {1{$random}};
  GEN_12 = GEN_76[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_77 = {1{$random}};
  GEN_13 = GEN_77[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_78 = {1{$random}};
  GEN_14 = GEN_78[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_79 = {1{$random}};
  GEN_15 = GEN_79[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_80 = {1{$random}};
  GEN_16 = GEN_80[11:0];
  `endif
  `ifdef RANDOMIZE
  GEN_81 = {2{$random}};
  GEN_17 = GEN_81[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_82 = {1{$random}};
  GEN_18 = GEN_82[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_83 = {1{$random}};
  GEN_19 = GEN_83[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_84 = {1{$random}};
  GEN_20 = GEN_84[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_85 = {1{$random}};
  GEN_21 = GEN_85[25:0];
  `endif
  `ifdef RANDOMIZE
  GEN_86 = {1{$random}};
  GEN_22 = GEN_86[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_87 = {1{$random}};
  GEN_23 = GEN_87[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_88 = {1{$random}};
  GEN_24 = GEN_88[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_89 = {2{$random}};
  GEN_25 = GEN_89[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_90 = {1{$random}};
  GEN_26 = GEN_90[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_91 = {1{$random}};
  GEN_27 = GEN_91[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_92 = {1{$random}};
  GEN_28 = GEN_92[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_93 = {1{$random}};
  GEN_29 = GEN_93[25:0];
  `endif
  `ifdef RANDOMIZE
  GEN_94 = {1{$random}};
  GEN_30 = GEN_94[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_95 = {1{$random}};
  GEN_31 = GEN_95[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_96 = {1{$random}};
  GEN_32 = GEN_96[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_97 = {2{$random}};
  GEN_33 = GEN_97[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_98 = {1{$random}};
  GEN_34 = GEN_98[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_99 = {1{$random}};
  GEN_35 = GEN_99[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_100 = {1{$random}};
  GEN_36 = GEN_100[25:0];
  `endif
  `ifdef RANDOMIZE
  GEN_101 = {1{$random}};
  GEN_37 = GEN_101[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_102 = {1{$random}};
  GEN_38 = GEN_102[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_103 = {1{$random}};
  GEN_39 = GEN_103[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_104 = {1{$random}};
  GEN_40 = GEN_104[25:0];
  `endif
  `ifdef RANDOMIZE
  GEN_105 = {1{$random}};
  GEN_41 = GEN_105[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_106 = {1{$random}};
  GEN_42 = GEN_106[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_107 = {1{$random}};
  GEN_43 = GEN_107[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_108 = {1{$random}};
  GEN_44 = GEN_108[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_109 = {1{$random}};
  GEN_45 = GEN_109[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_110 = {1{$random}};
  GEN_46 = GEN_110[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_111 = {1{$random}};
  GEN_47 = GEN_111[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_112 = {1{$random}};
  GEN_48 = GEN_112[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_113 = {2{$random}};
  GEN_49 = GEN_113[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_114 = {1{$random}};
  GEN_50 = GEN_114[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_115 = {1{$random}};
  GEN_51 = GEN_115[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_116 = {1{$random}};
  GEN_52 = GEN_116[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_117 = {1{$random}};
  GEN_53 = GEN_117[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_118 = {1{$random}};
  GEN_54 = GEN_118[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_119 = {1{$random}};
  GEN_55 = GEN_119[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_120 = {1{$random}};
  GEN_56 = GEN_120[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_121 = {2{$random}};
  GEN_57 = GEN_121[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_122 = {1{$random}};
  GEN_58 = GEN_122[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_123 = {1{$random}};
  GEN_59 = GEN_123[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_124 = {1{$random}};
  GEN_60 = GEN_124[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_125 = {1{$random}};
  GEN_61 = GEN_125[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_126 = {1{$random}};
  GEN_62 = GEN_126[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_127 = {1{$random}};
  GEN_63 = GEN_127[1:0];
  `endif
  end
`endif
endmodule
module ManagerToClientStatelessBridge(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input   io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [11:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output  io_inner_grant_bits_client_xact_id,
  output [1:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [1:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input   io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [1:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [11:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [1:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [1:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id
);
  wire [1:0] T_1215;
  wire [1:0] T_1216;
  wire  T_1217;
  wire  T_1218;
  wire  T_1224;
  wire  T_1225;
  wire  T_1227;
  reg [25:0] GEN_0;
  reg [31:0] GEN_5;
  reg [1:0] GEN_1;
  reg [31:0] GEN_6;
  reg  GEN_2;
  reg [31:0] GEN_7;
  reg  GEN_3;
  reg [31:0] GEN_8;
  reg  GEN_4;
  reg [31:0] GEN_9;
  assign io_inner_acquire_ready = io_outer_acquire_ready;
  assign io_inner_grant_valid = io_outer_grant_valid;
  assign io_inner_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign io_inner_grant_bits_client_xact_id = T_1217;
  assign io_inner_grant_bits_manager_xact_id = {{1'd0}, io_outer_grant_bits_manager_xact_id};
  assign io_inner_grant_bits_is_builtin_type = io_outer_grant_bits_is_builtin_type;
  assign io_inner_grant_bits_g_type = io_outer_grant_bits_g_type;
  assign io_inner_grant_bits_data = io_outer_grant_bits_data;
  assign io_inner_grant_bits_client_id = T_1218;
  assign io_inner_finish_ready = 1'h1;
  assign io_inner_probe_valid = 1'h0;
  assign io_inner_probe_bits_addr_block = GEN_0;
  assign io_inner_probe_bits_p_type = GEN_1;
  assign io_inner_probe_bits_client_id = GEN_2;
  assign io_inner_release_ready = io_outer_release_ready;
  assign io_outer_acquire_valid = io_inner_acquire_valid;
  assign io_outer_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign io_outer_acquire_bits_client_xact_id = T_1215;
  assign io_outer_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign io_outer_acquire_bits_union = io_inner_acquire_bits_union;
  assign io_outer_acquire_bits_data = io_inner_acquire_bits_data;
  assign io_outer_probe_ready = 1'h0;
  assign io_outer_release_valid = io_inner_release_valid;
  assign io_outer_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_release_bits_client_xact_id = T_1216;
  assign io_outer_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign io_outer_release_bits_r_type = io_inner_release_bits_r_type;
  assign io_outer_release_bits_data = io_inner_release_bits_data;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_finish_valid = 1'h0;
  assign io_outer_finish_bits_manager_xact_id = GEN_3;
  assign io_outer_finish_bits_manager_id = GEN_4;
  assign T_1215 = {io_inner_acquire_bits_client_id,io_inner_acquire_bits_client_xact_id};
  assign T_1216 = {io_inner_release_bits_client_id,io_inner_release_bits_client_xact_id};
  assign T_1217 = io_outer_grant_bits_client_xact_id[0];
  assign T_1218 = io_outer_grant_bits_client_xact_id[1];
  assign T_1224 = io_outer_probe_valid == 1'h0;
  assign T_1225 = T_1224 | reset;
  assign T_1227 = T_1225 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_5 = {1{$random}};
  GEN_0 = GEN_5[25:0];
  `endif
  `ifdef RANDOMIZE
  GEN_6 = {1{$random}};
  GEN_1 = GEN_6[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_7 = {1{$random}};
  GEN_2 = GEN_7[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_8 = {1{$random}};
  GEN_3 = GEN_8[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_9 = {1{$random}};
  GEN_4 = GEN_9[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1227) begin
          $fwrite(32'h80000002,"Assertion failed: L2 agent got illegal probe\n    at Agents.scala:159 assert(!io.outer.probe.valid, ---L2 agent got illegal probe---)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1227) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module MMIOTileLinkManager(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input   io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [11:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output  io_inner_grant_bits_client_xact_id,
  output [1:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [1:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input   io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [1:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [11:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [1:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data
);
  wire  T_880;
  wire [2:0] T_889_0;
  wire  T_891;
  wire  T_892;
  wire  multibeat_fire;
  wire  T_894;
  wire  multibeat_start;
  wire  T_896;
  wire  multibeat_end;
  reg [3:0] xact_pending;
  reg [31:0] GEN_33;
  wire [3:0] T_898;
  wire  T_899;
  wire  T_900;
  wire  T_901;
  wire [1:0] T_907;
  wire [1:0] T_908;
  wire [1:0] xact_id_sel;
  reg [1:0] xact_id_reg;
  reg [31:0] GEN_34;
  wire [1:0] GEN_4;
  reg  xact_multibeat;
  reg [31:0] GEN_35;
  wire [1:0] outer_xact_id;
  wire  T_912;
  wire  xact_free;
  reg  xact_buffer_0_client_id;
  reg [31:0] GEN_36;
  reg  xact_buffer_0_client_xact_id;
  reg [31:0] GEN_37;
  reg  xact_buffer_1_client_id;
  reg [31:0] GEN_38;
  reg  xact_buffer_1_client_xact_id;
  reg [31:0] GEN_39;
  reg  xact_buffer_2_client_id;
  reg [31:0] GEN_40;
  reg  xact_buffer_2_client_xact_id;
  reg [31:0] GEN_41;
  reg  xact_buffer_3_client_id;
  reg [31:0] GEN_42;
  reg  xact_buffer_3_client_xact_id;
  reg [31:0] GEN_43;
  wire  T_1229;
  wire  T_1230;
  wire [2:0] T_1240_0;
  wire  T_1242;
  wire  T_1243;
  wire  T_1245;
  wire  T_1248;
  wire  T_1249;
  wire [3:0] T_1251;
  wire [3:0] T_1253;
  wire [3:0] T_1254;
  wire  T_1255;
  wire [3:0] T_1257;
  wire [3:0] T_1259;
  wire [3:0] T_1260;
  wire [3:0] T_1261;
  wire  T_1262;
  wire [2:0] T_1270_0;
  wire [3:0] GEN_31;
  wire  T_1272;
  wire  T_1273;
  wire  T_1274;
  wire  T_1277;
  wire  T_1279;
  wire  T_1280;
  wire  T_1281;
  wire  T_1287;
  wire  T_1289;
  wire  T_1292;
  wire  T_1293;
  wire [3:0] T_1295;
  wire [3:0] T_1297;
  wire [3:0] T_1298;
  wire [3:0] T_1299;
  wire [2:0] T_1309_0;
  wire  T_1311;
  wire  T_1312;
  wire  T_1314;
  wire  T_1317;
  wire  T_1318;
  wire  GEN_0;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_1;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire  GEN_17;
  wire  GEN_19;
  wire  GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire  GEN_2;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire  GEN_3;
  wire  GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  reg [25:0] GEN_13;
  reg [31:0] GEN_44;
  reg [1:0] GEN_18;
  reg [31:0] GEN_45;
  reg  GEN_32;
  reg [31:0] GEN_46;
  assign io_inner_acquire_ready = T_1229;
  assign io_inner_grant_valid = io_outer_grant_valid;
  assign io_inner_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign io_inner_grant_bits_client_xact_id = GEN_3;
  assign io_inner_grant_bits_manager_xact_id = io_outer_grant_bits_client_xact_id;
  assign io_inner_grant_bits_is_builtin_type = io_outer_grant_bits_is_builtin_type;
  assign io_inner_grant_bits_g_type = io_outer_grant_bits_g_type;
  assign io_inner_grant_bits_data = io_outer_grant_bits_data;
  assign io_inner_grant_bits_client_id = GEN_2;
  assign io_inner_finish_ready = 1'h1;
  assign io_inner_probe_valid = 1'h0;
  assign io_inner_probe_bits_addr_block = GEN_13;
  assign io_inner_probe_bits_p_type = GEN_18;
  assign io_inner_probe_bits_client_id = GEN_32;
  assign io_inner_release_ready = 1'h0;
  assign io_outer_acquire_valid = T_1230;
  assign io_outer_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign io_outer_acquire_bits_client_xact_id = outer_xact_id;
  assign io_outer_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign io_outer_acquire_bits_union = io_inner_acquire_bits_union;
  assign io_outer_acquire_bits_data = io_inner_acquire_bits_data;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign T_880 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T_889_0 = 3'h3;
  assign T_891 = io_outer_acquire_bits_a_type == T_889_0;
  assign T_892 = io_outer_acquire_bits_is_builtin_type & T_891;
  assign multibeat_fire = T_880 & T_892;
  assign T_894 = io_outer_acquire_bits_addr_beat == 3'h0;
  assign multibeat_start = multibeat_fire & T_894;
  assign T_896 = io_outer_acquire_bits_addr_beat == 3'h7;
  assign multibeat_end = multibeat_fire & T_896;
  assign T_898 = ~ xact_pending;
  assign T_899 = T_898[0];
  assign T_900 = T_898[1];
  assign T_901 = T_898[2];
  assign T_907 = T_901 ? 2'h2 : 2'h3;
  assign T_908 = T_900 ? 2'h1 : T_907;
  assign xact_id_sel = T_899 ? 2'h0 : T_908;
  assign GEN_4 = multibeat_start ? xact_id_sel : xact_id_reg;
  assign outer_xact_id = xact_multibeat ? xact_id_reg : xact_id_sel;
  assign T_912 = T_898 == 4'h0;
  assign xact_free = T_912 == 1'h0;
  assign T_1229 = io_outer_acquire_ready & xact_free;
  assign T_1230 = io_inner_acquire_valid & xact_free;
  assign T_1240_0 = 3'h3;
  assign T_1242 = io_outer_acquire_bits_a_type == T_1240_0;
  assign T_1243 = io_outer_acquire_bits_is_builtin_type & T_1242;
  assign T_1245 = T_1243 == 1'h0;
  assign T_1248 = T_1245 | T_896;
  assign T_1249 = T_880 & T_1248;
  assign T_1251 = 4'h1 << io_outer_acquire_bits_client_xact_id;
  assign T_1253 = T_1249 ? T_1251 : 4'h0;
  assign T_1254 = xact_pending | T_1253;
  assign T_1255 = io_inner_finish_ready & io_inner_finish_valid;
  assign T_1257 = 4'h1 << io_inner_finish_bits_manager_xact_id;
  assign T_1259 = T_1255 ? T_1257 : 4'h0;
  assign T_1260 = ~ T_1259;
  assign T_1261 = T_1254 & T_1260;
  assign T_1262 = io_inner_grant_ready & io_inner_grant_valid;
  assign T_1270_0 = 3'h5;
  assign GEN_31 = {{1'd0}, T_1270_0};
  assign T_1272 = io_inner_grant_bits_g_type == GEN_31;
  assign T_1273 = io_inner_grant_bits_g_type == 4'h0;
  assign T_1274 = io_inner_grant_bits_is_builtin_type ? T_1272 : T_1273;
  assign T_1277 = T_1274 == 1'h0;
  assign T_1279 = io_inner_grant_bits_addr_beat == 3'h7;
  assign T_1280 = T_1277 | T_1279;
  assign T_1281 = T_1262 & T_1280;
  assign T_1287 = io_inner_grant_bits_is_builtin_type & T_1273;
  assign T_1289 = T_1287 == 1'h0;
  assign T_1292 = T_1289 == 1'h0;
  assign T_1293 = T_1281 & T_1292;
  assign T_1295 = 4'h1 << io_inner_grant_bits_manager_xact_id;
  assign T_1297 = T_1293 ? T_1295 : 4'h0;
  assign T_1298 = ~ T_1297;
  assign T_1299 = T_1261 & T_1298;
  assign T_1309_0 = 3'h3;
  assign T_1311 = io_outer_acquire_bits_a_type == T_1309_0;
  assign T_1312 = io_outer_acquire_bits_is_builtin_type & T_1311;
  assign T_1314 = T_1312 == 1'h0;
  assign T_1317 = T_1314 | T_896;
  assign T_1318 = T_880 & T_1317;
  assign GEN_0 = io_inner_acquire_bits_client_id;
  assign GEN_5 = 2'h0 == outer_xact_id ? GEN_0 : xact_buffer_0_client_id;
  assign GEN_6 = 2'h1 == outer_xact_id ? GEN_0 : xact_buffer_1_client_id;
  assign GEN_7 = 2'h2 == outer_xact_id ? GEN_0 : xact_buffer_2_client_id;
  assign GEN_8 = 2'h3 == outer_xact_id ? GEN_0 : xact_buffer_3_client_id;
  assign GEN_1 = io_inner_acquire_bits_client_xact_id;
  assign GEN_9 = 2'h0 == outer_xact_id ? GEN_1 : xact_buffer_0_client_xact_id;
  assign GEN_10 = 2'h1 == outer_xact_id ? GEN_1 : xact_buffer_1_client_xact_id;
  assign GEN_11 = 2'h2 == outer_xact_id ? GEN_1 : xact_buffer_2_client_xact_id;
  assign GEN_12 = 2'h3 == outer_xact_id ? GEN_1 : xact_buffer_3_client_xact_id;
  assign GEN_14 = T_1318 ? GEN_5 : xact_buffer_0_client_id;
  assign GEN_15 = T_1318 ? GEN_6 : xact_buffer_1_client_id;
  assign GEN_16 = T_1318 ? GEN_7 : xact_buffer_2_client_id;
  assign GEN_17 = T_1318 ? GEN_8 : xact_buffer_3_client_id;
  assign GEN_19 = T_1318 ? GEN_9 : xact_buffer_0_client_xact_id;
  assign GEN_20 = T_1318 ? GEN_10 : xact_buffer_1_client_xact_id;
  assign GEN_21 = T_1318 ? GEN_11 : xact_buffer_2_client_xact_id;
  assign GEN_22 = T_1318 ? GEN_12 : xact_buffer_3_client_xact_id;
  assign GEN_23 = multibeat_start ? 1'h1 : xact_multibeat;
  assign GEN_24 = multibeat_end ? 1'h0 : GEN_23;
  assign GEN_2 = GEN_27;
  assign GEN_25 = 2'h1 == io_outer_grant_bits_client_xact_id ? xact_buffer_1_client_id : xact_buffer_0_client_id;
  assign GEN_26 = 2'h2 == io_outer_grant_bits_client_xact_id ? xact_buffer_2_client_id : GEN_25;
  assign GEN_27 = 2'h3 == io_outer_grant_bits_client_xact_id ? xact_buffer_3_client_id : GEN_26;
  assign GEN_3 = GEN_30;
  assign GEN_28 = 2'h1 == io_outer_grant_bits_client_xact_id ? xact_buffer_1_client_xact_id : xact_buffer_0_client_xact_id;
  assign GEN_29 = 2'h2 == io_outer_grant_bits_client_xact_id ? xact_buffer_2_client_xact_id : GEN_28;
  assign GEN_30 = 2'h3 == io_outer_grant_bits_client_xact_id ? xact_buffer_3_client_xact_id : GEN_29;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_33 = {1{$random}};
  xact_pending = GEN_33[3:0];
  `endif
  `ifdef RANDOMIZE
  GEN_34 = {1{$random}};
  xact_id_reg = GEN_34[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_35 = {1{$random}};
  xact_multibeat = GEN_35[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_36 = {1{$random}};
  xact_buffer_0_client_id = GEN_36[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_37 = {1{$random}};
  xact_buffer_0_client_xact_id = GEN_37[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_38 = {1{$random}};
  xact_buffer_1_client_id = GEN_38[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_39 = {1{$random}};
  xact_buffer_1_client_xact_id = GEN_39[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_40 = {1{$random}};
  xact_buffer_2_client_id = GEN_40[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_41 = {1{$random}};
  xact_buffer_2_client_xact_id = GEN_41[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_42 = {1{$random}};
  xact_buffer_3_client_id = GEN_42[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_43 = {1{$random}};
  xact_buffer_3_client_xact_id = GEN_43[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_44 = {1{$random}};
  GEN_13 = GEN_44[25:0];
  `endif
  `ifdef RANDOMIZE
  GEN_45 = {1{$random}};
  GEN_18 = GEN_45[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_46 = {1{$random}};
  GEN_32 = GEN_46[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      xact_pending <= 4'h0;
    end else begin
      xact_pending <= T_1299;
    end
    if(1'h0) begin
    end else begin
      if(multibeat_start) begin
        if(T_899) begin
          xact_id_reg <= 2'h0;
        end else begin
          if(T_900) begin
            xact_id_reg <= 2'h1;
          end else begin
            if(T_901) begin
              xact_id_reg <= 2'h2;
            end else begin
              xact_id_reg <= 2'h3;
            end
          end
        end
      end
    end
    if(reset) begin
      xact_multibeat <= 1'h0;
    end else begin
      if(multibeat_end) begin
        xact_multibeat <= 1'h0;
      end else begin
        if(multibeat_start) begin
          xact_multibeat <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1318) begin
        if(2'h0 == outer_xact_id) begin
          xact_buffer_0_client_id <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1318) begin
        if(2'h0 == outer_xact_id) begin
          xact_buffer_0_client_xact_id <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1318) begin
        if(2'h1 == outer_xact_id) begin
          xact_buffer_1_client_id <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1318) begin
        if(2'h1 == outer_xact_id) begin
          xact_buffer_1_client_xact_id <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1318) begin
        if(2'h2 == outer_xact_id) begin
          xact_buffer_2_client_id <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1318) begin
        if(2'h2 == outer_xact_id) begin
          xact_buffer_2_client_xact_id <= GEN_1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1318) begin
        if(2'h3 == outer_xact_id) begin
          xact_buffer_3_client_id <= GEN_0;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1318) begin
        if(2'h3 == outer_xact_id) begin
          xact_buffer_3_client_xact_id <= GEN_1;
        end
      end
    end
  end
endmodule
module Queue_8(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [25:0] io_enq_bits_addr_block,
  input  [1:0] io_enq_bits_client_xact_id,
  input  [2:0] io_enq_bits_addr_beat,
  input   io_enq_bits_is_builtin_type,
  input  [2:0] io_enq_bits_a_type,
  input  [11:0] io_enq_bits_union,
  input  [63:0] io_enq_bits_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [25:0] io_deq_bits_addr_block,
  output [1:0] io_deq_bits_client_xact_id,
  output [2:0] io_deq_bits_addr_beat,
  output  io_deq_bits_is_builtin_type,
  output [2:0] io_deq_bits_a_type,
  output [11:0] io_deq_bits_union,
  output [63:0] io_deq_bits_data,
  output  io_count
);
  reg [25:0] ram_addr_block [0:0];
  reg [31:0] GEN_0;
  wire [25:0] ram_addr_block_T_254_data;
  wire  ram_addr_block_T_254_addr;
  wire  ram_addr_block_T_254_en;
  wire [25:0] ram_addr_block_T_224_data;
  wire  ram_addr_block_T_224_addr;
  wire  ram_addr_block_T_224_mask;
  wire  ram_addr_block_T_224_en;
  reg [1:0] ram_client_xact_id [0:0];
  reg [31:0] GEN_1;
  wire [1:0] ram_client_xact_id_T_254_data;
  wire  ram_client_xact_id_T_254_addr;
  wire  ram_client_xact_id_T_254_en;
  wire [1:0] ram_client_xact_id_T_224_data;
  wire  ram_client_xact_id_T_224_addr;
  wire  ram_client_xact_id_T_224_mask;
  wire  ram_client_xact_id_T_224_en;
  reg [2:0] ram_addr_beat [0:0];
  reg [31:0] GEN_2;
  wire [2:0] ram_addr_beat_T_254_data;
  wire  ram_addr_beat_T_254_addr;
  wire  ram_addr_beat_T_254_en;
  wire [2:0] ram_addr_beat_T_224_data;
  wire  ram_addr_beat_T_224_addr;
  wire  ram_addr_beat_T_224_mask;
  wire  ram_addr_beat_T_224_en;
  reg  ram_is_builtin_type [0:0];
  reg [31:0] GEN_3;
  wire  ram_is_builtin_type_T_254_data;
  wire  ram_is_builtin_type_T_254_addr;
  wire  ram_is_builtin_type_T_254_en;
  wire  ram_is_builtin_type_T_224_data;
  wire  ram_is_builtin_type_T_224_addr;
  wire  ram_is_builtin_type_T_224_mask;
  wire  ram_is_builtin_type_T_224_en;
  reg [2:0] ram_a_type [0:0];
  reg [31:0] GEN_4;
  wire [2:0] ram_a_type_T_254_data;
  wire  ram_a_type_T_254_addr;
  wire  ram_a_type_T_254_en;
  wire [2:0] ram_a_type_T_224_data;
  wire  ram_a_type_T_224_addr;
  wire  ram_a_type_T_224_mask;
  wire  ram_a_type_T_224_en;
  reg [11:0] ram_union [0:0];
  reg [31:0] GEN_5;
  wire [11:0] ram_union_T_254_data;
  wire  ram_union_T_254_addr;
  wire  ram_union_T_254_en;
  wire [11:0] ram_union_T_224_data;
  wire  ram_union_T_224_addr;
  wire  ram_union_T_224_mask;
  wire  ram_union_T_224_en;
  reg [63:0] ram_data [0:0];
  reg [63:0] GEN_6;
  wire [63:0] ram_data_T_254_data;
  wire  ram_data_T_254_addr;
  wire  ram_data_T_254_en;
  wire [63:0] ram_data_T_224_data;
  wire  ram_data_T_224_addr;
  wire  ram_data_T_224_mask;
  wire  ram_data_T_224_en;
  reg  maybe_full;
  reg [31:0] GEN_7;
  wire  T_221;
  wire  T_222;
  wire  do_enq;
  wire  T_223;
  wire  do_deq;
  wire  T_249;
  wire  GEN_17;
  wire  T_251;
  wire [1:0] T_277;
  wire  ptr_diff;
  wire [1:0] T_279;
  assign io_enq_ready = T_221;
  assign io_deq_valid = T_251;
  assign io_deq_bits_addr_block = ram_addr_block_T_254_data;
  assign io_deq_bits_client_xact_id = ram_client_xact_id_T_254_data;
  assign io_deq_bits_addr_beat = ram_addr_beat_T_254_data;
  assign io_deq_bits_is_builtin_type = ram_is_builtin_type_T_254_data;
  assign io_deq_bits_a_type = ram_a_type_T_254_data;
  assign io_deq_bits_union = ram_union_T_254_data;
  assign io_deq_bits_data = ram_data_T_254_data;
  assign io_count = T_279[0];
  assign ram_addr_block_T_254_addr = 1'h0;
  assign ram_addr_block_T_254_en = 1'h1;
  assign ram_addr_block_T_254_data = ram_addr_block[ram_addr_block_T_254_addr];
  assign ram_addr_block_T_224_data = io_enq_bits_addr_block;
  assign ram_addr_block_T_224_addr = 1'h0;
  assign ram_addr_block_T_224_mask = do_enq;
  assign ram_addr_block_T_224_en = do_enq;
  assign ram_client_xact_id_T_254_addr = 1'h0;
  assign ram_client_xact_id_T_254_en = 1'h1;
  assign ram_client_xact_id_T_254_data = ram_client_xact_id[ram_client_xact_id_T_254_addr];
  assign ram_client_xact_id_T_224_data = io_enq_bits_client_xact_id;
  assign ram_client_xact_id_T_224_addr = 1'h0;
  assign ram_client_xact_id_T_224_mask = do_enq;
  assign ram_client_xact_id_T_224_en = do_enq;
  assign ram_addr_beat_T_254_addr = 1'h0;
  assign ram_addr_beat_T_254_en = 1'h1;
  assign ram_addr_beat_T_254_data = ram_addr_beat[ram_addr_beat_T_254_addr];
  assign ram_addr_beat_T_224_data = io_enq_bits_addr_beat;
  assign ram_addr_beat_T_224_addr = 1'h0;
  assign ram_addr_beat_T_224_mask = do_enq;
  assign ram_addr_beat_T_224_en = do_enq;
  assign ram_is_builtin_type_T_254_addr = 1'h0;
  assign ram_is_builtin_type_T_254_en = 1'h1;
  assign ram_is_builtin_type_T_254_data = ram_is_builtin_type[ram_is_builtin_type_T_254_addr];
  assign ram_is_builtin_type_T_224_data = io_enq_bits_is_builtin_type;
  assign ram_is_builtin_type_T_224_addr = 1'h0;
  assign ram_is_builtin_type_T_224_mask = do_enq;
  assign ram_is_builtin_type_T_224_en = do_enq;
  assign ram_a_type_T_254_addr = 1'h0;
  assign ram_a_type_T_254_en = 1'h1;
  assign ram_a_type_T_254_data = ram_a_type[ram_a_type_T_254_addr];
  assign ram_a_type_T_224_data = io_enq_bits_a_type;
  assign ram_a_type_T_224_addr = 1'h0;
  assign ram_a_type_T_224_mask = do_enq;
  assign ram_a_type_T_224_en = do_enq;
  assign ram_union_T_254_addr = 1'h0;
  assign ram_union_T_254_en = 1'h1;
  assign ram_union_T_254_data = ram_union[ram_union_T_254_addr];
  assign ram_union_T_224_data = io_enq_bits_union;
  assign ram_union_T_224_addr = 1'h0;
  assign ram_union_T_224_mask = do_enq;
  assign ram_union_T_224_en = do_enq;
  assign ram_data_T_254_addr = 1'h0;
  assign ram_data_T_254_en = 1'h1;
  assign ram_data_T_254_data = ram_data[ram_data_T_254_addr];
  assign ram_data_T_224_data = io_enq_bits_data;
  assign ram_data_T_224_addr = 1'h0;
  assign ram_data_T_224_mask = do_enq;
  assign ram_data_T_224_en = do_enq;
  assign T_221 = maybe_full == 1'h0;
  assign T_222 = io_enq_ready & io_enq_valid;
  assign do_enq = T_222;
  assign T_223 = io_deq_ready & io_deq_valid;
  assign do_deq = T_223;
  assign T_249 = do_enq != do_deq;
  assign GEN_17 = T_249 ? do_enq : maybe_full;
  assign T_251 = T_221 == 1'h0;
  assign T_277 = 1'h0 - 1'h0;
  assign ptr_diff = T_277[0:0];
  assign T_279 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr_block[initvar] = GEN_0[25:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_client_xact_id[initvar] = GEN_1[1:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr_beat[initvar] = GEN_2[2:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_is_builtin_type[initvar] = GEN_3[0:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_a_type[initvar] = GEN_4[2:0];
  `endif
  GEN_5 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_union[initvar] = GEN_5[11:0];
  `endif
  GEN_6 = {2{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = GEN_6[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_7 = {1{$random}};
  maybe_full = GEN_7[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_addr_block_T_224_en & ram_addr_block_T_224_mask) begin
      ram_addr_block[ram_addr_block_T_224_addr] <= ram_addr_block_T_224_data;
    end
    if(ram_client_xact_id_T_224_en & ram_client_xact_id_T_224_mask) begin
      ram_client_xact_id[ram_client_xact_id_T_224_addr] <= ram_client_xact_id_T_224_data;
    end
    if(ram_addr_beat_T_224_en & ram_addr_beat_T_224_mask) begin
      ram_addr_beat[ram_addr_beat_T_224_addr] <= ram_addr_beat_T_224_data;
    end
    if(ram_is_builtin_type_T_224_en & ram_is_builtin_type_T_224_mask) begin
      ram_is_builtin_type[ram_is_builtin_type_T_224_addr] <= ram_is_builtin_type_T_224_data;
    end
    if(ram_a_type_T_224_en & ram_a_type_T_224_mask) begin
      ram_a_type[ram_a_type_T_224_addr] <= ram_a_type_T_224_data;
    end
    if(ram_union_T_224_en & ram_union_T_224_mask) begin
      ram_union[ram_union_T_224_addr] <= ram_union_T_224_data;
    end
    if(ram_data_T_224_en & ram_data_T_224_mask) begin
      ram_data[ram_data_T_224_addr] <= ram_data_T_224_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_249) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_9(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [2:0] io_enq_bits_addr_beat,
  input  [1:0] io_enq_bits_client_xact_id,
  input   io_enq_bits_manager_xact_id,
  input   io_enq_bits_is_builtin_type,
  input  [3:0] io_enq_bits_g_type,
  input  [63:0] io_enq_bits_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [2:0] io_deq_bits_addr_beat,
  output [1:0] io_deq_bits_client_xact_id,
  output  io_deq_bits_manager_xact_id,
  output  io_deq_bits_is_builtin_type,
  output [3:0] io_deq_bits_g_type,
  output [63:0] io_deq_bits_data,
  output  io_count
);
  reg [2:0] ram_addr_beat [0:0];
  reg [31:0] GEN_0;
  wire [2:0] ram_addr_beat_T_244_data;
  wire  ram_addr_beat_T_244_addr;
  wire  ram_addr_beat_T_244_en;
  wire [2:0] ram_addr_beat_T_215_data;
  wire  ram_addr_beat_T_215_addr;
  wire  ram_addr_beat_T_215_mask;
  wire  ram_addr_beat_T_215_en;
  reg [1:0] ram_client_xact_id [0:0];
  reg [31:0] GEN_1;
  wire [1:0] ram_client_xact_id_T_244_data;
  wire  ram_client_xact_id_T_244_addr;
  wire  ram_client_xact_id_T_244_en;
  wire [1:0] ram_client_xact_id_T_215_data;
  wire  ram_client_xact_id_T_215_addr;
  wire  ram_client_xact_id_T_215_mask;
  wire  ram_client_xact_id_T_215_en;
  reg  ram_manager_xact_id [0:0];
  reg [31:0] GEN_2;
  wire  ram_manager_xact_id_T_244_data;
  wire  ram_manager_xact_id_T_244_addr;
  wire  ram_manager_xact_id_T_244_en;
  wire  ram_manager_xact_id_T_215_data;
  wire  ram_manager_xact_id_T_215_addr;
  wire  ram_manager_xact_id_T_215_mask;
  wire  ram_manager_xact_id_T_215_en;
  reg  ram_is_builtin_type [0:0];
  reg [31:0] GEN_3;
  wire  ram_is_builtin_type_T_244_data;
  wire  ram_is_builtin_type_T_244_addr;
  wire  ram_is_builtin_type_T_244_en;
  wire  ram_is_builtin_type_T_215_data;
  wire  ram_is_builtin_type_T_215_addr;
  wire  ram_is_builtin_type_T_215_mask;
  wire  ram_is_builtin_type_T_215_en;
  reg [3:0] ram_g_type [0:0];
  reg [31:0] GEN_4;
  wire [3:0] ram_g_type_T_244_data;
  wire  ram_g_type_T_244_addr;
  wire  ram_g_type_T_244_en;
  wire [3:0] ram_g_type_T_215_data;
  wire  ram_g_type_T_215_addr;
  wire  ram_g_type_T_215_mask;
  wire  ram_g_type_T_215_en;
  reg [63:0] ram_data [0:0];
  reg [63:0] GEN_5;
  wire [63:0] ram_data_T_244_data;
  wire  ram_data_T_244_addr;
  wire  ram_data_T_244_en;
  wire [63:0] ram_data_T_215_data;
  wire  ram_data_T_215_addr;
  wire  ram_data_T_215_mask;
  wire  ram_data_T_215_en;
  reg  maybe_full;
  reg [31:0] GEN_6;
  wire  T_212;
  wire  T_213;
  wire  do_enq;
  wire  T_214;
  wire  do_deq;
  wire  T_239;
  wire  GEN_15;
  wire  T_241;
  wire [1:0] T_266;
  wire  ptr_diff;
  wire [1:0] T_268;
  assign io_enq_ready = T_212;
  assign io_deq_valid = T_241;
  assign io_deq_bits_addr_beat = ram_addr_beat_T_244_data;
  assign io_deq_bits_client_xact_id = ram_client_xact_id_T_244_data;
  assign io_deq_bits_manager_xact_id = ram_manager_xact_id_T_244_data;
  assign io_deq_bits_is_builtin_type = ram_is_builtin_type_T_244_data;
  assign io_deq_bits_g_type = ram_g_type_T_244_data;
  assign io_deq_bits_data = ram_data_T_244_data;
  assign io_count = T_268[0];
  assign ram_addr_beat_T_244_addr = 1'h0;
  assign ram_addr_beat_T_244_en = 1'h1;
  assign ram_addr_beat_T_244_data = ram_addr_beat[ram_addr_beat_T_244_addr];
  assign ram_addr_beat_T_215_data = io_enq_bits_addr_beat;
  assign ram_addr_beat_T_215_addr = 1'h0;
  assign ram_addr_beat_T_215_mask = do_enq;
  assign ram_addr_beat_T_215_en = do_enq;
  assign ram_client_xact_id_T_244_addr = 1'h0;
  assign ram_client_xact_id_T_244_en = 1'h1;
  assign ram_client_xact_id_T_244_data = ram_client_xact_id[ram_client_xact_id_T_244_addr];
  assign ram_client_xact_id_T_215_data = io_enq_bits_client_xact_id;
  assign ram_client_xact_id_T_215_addr = 1'h0;
  assign ram_client_xact_id_T_215_mask = do_enq;
  assign ram_client_xact_id_T_215_en = do_enq;
  assign ram_manager_xact_id_T_244_addr = 1'h0;
  assign ram_manager_xact_id_T_244_en = 1'h1;
  assign ram_manager_xact_id_T_244_data = ram_manager_xact_id[ram_manager_xact_id_T_244_addr];
  assign ram_manager_xact_id_T_215_data = io_enq_bits_manager_xact_id;
  assign ram_manager_xact_id_T_215_addr = 1'h0;
  assign ram_manager_xact_id_T_215_mask = do_enq;
  assign ram_manager_xact_id_T_215_en = do_enq;
  assign ram_is_builtin_type_T_244_addr = 1'h0;
  assign ram_is_builtin_type_T_244_en = 1'h1;
  assign ram_is_builtin_type_T_244_data = ram_is_builtin_type[ram_is_builtin_type_T_244_addr];
  assign ram_is_builtin_type_T_215_data = io_enq_bits_is_builtin_type;
  assign ram_is_builtin_type_T_215_addr = 1'h0;
  assign ram_is_builtin_type_T_215_mask = do_enq;
  assign ram_is_builtin_type_T_215_en = do_enq;
  assign ram_g_type_T_244_addr = 1'h0;
  assign ram_g_type_T_244_en = 1'h1;
  assign ram_g_type_T_244_data = ram_g_type[ram_g_type_T_244_addr];
  assign ram_g_type_T_215_data = io_enq_bits_g_type;
  assign ram_g_type_T_215_addr = 1'h0;
  assign ram_g_type_T_215_mask = do_enq;
  assign ram_g_type_T_215_en = do_enq;
  assign ram_data_T_244_addr = 1'h0;
  assign ram_data_T_244_en = 1'h1;
  assign ram_data_T_244_data = ram_data[ram_data_T_244_addr];
  assign ram_data_T_215_data = io_enq_bits_data;
  assign ram_data_T_215_addr = 1'h0;
  assign ram_data_T_215_mask = do_enq;
  assign ram_data_T_215_en = do_enq;
  assign T_212 = maybe_full == 1'h0;
  assign T_213 = io_enq_ready & io_enq_valid;
  assign do_enq = T_213;
  assign T_214 = io_deq_ready & io_deq_valid;
  assign do_deq = T_214;
  assign T_239 = do_enq != do_deq;
  assign GEN_15 = T_239 ? do_enq : maybe_full;
  assign T_241 = T_212 == 1'h0;
  assign T_266 = 1'h0 - 1'h0;
  assign ptr_diff = T_266[0:0];
  assign T_268 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr_beat[initvar] = GEN_0[2:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_client_xact_id[initvar] = GEN_1[1:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_manager_xact_id[initvar] = GEN_2[0:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_is_builtin_type[initvar] = GEN_3[0:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_g_type[initvar] = GEN_4[3:0];
  `endif
  GEN_5 = {2{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = GEN_5[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_6 = {1{$random}};
  maybe_full = GEN_6[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_addr_beat_T_215_en & ram_addr_beat_T_215_mask) begin
      ram_addr_beat[ram_addr_beat_T_215_addr] <= ram_addr_beat_T_215_data;
    end
    if(ram_client_xact_id_T_215_en & ram_client_xact_id_T_215_mask) begin
      ram_client_xact_id[ram_client_xact_id_T_215_addr] <= ram_client_xact_id_T_215_data;
    end
    if(ram_manager_xact_id_T_215_en & ram_manager_xact_id_T_215_mask) begin
      ram_manager_xact_id[ram_manager_xact_id_T_215_addr] <= ram_manager_xact_id_T_215_data;
    end
    if(ram_is_builtin_type_T_215_en & ram_is_builtin_type_T_215_mask) begin
      ram_is_builtin_type[ram_is_builtin_type_T_215_addr] <= ram_is_builtin_type_T_215_data;
    end
    if(ram_g_type_T_215_en & ram_g_type_T_215_mask) begin
      ram_g_type[ram_g_type_T_215_addr] <= ram_g_type_T_215_data;
    end
    if(ram_data_T_215_en & ram_data_T_215_mask) begin
      ram_data[ram_data_T_215_addr] <= ram_data_T_215_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_239) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module ClientUncachedTileLinkIOArbiter_1(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_acquire_ready,
  output  io_out_acquire_valid,
  output [25:0] io_out_acquire_bits_addr_block,
  output [1:0] io_out_acquire_bits_client_xact_id,
  output [2:0] io_out_acquire_bits_addr_beat,
  output  io_out_acquire_bits_is_builtin_type,
  output [2:0] io_out_acquire_bits_a_type,
  output [11:0] io_out_acquire_bits_union,
  output [63:0] io_out_acquire_bits_data,
  output  io_out_grant_ready,
  input   io_out_grant_valid,
  input  [2:0] io_out_grant_bits_addr_beat,
  input  [1:0] io_out_grant_bits_client_xact_id,
  input   io_out_grant_bits_manager_xact_id,
  input   io_out_grant_bits_is_builtin_type,
  input  [3:0] io_out_grant_bits_g_type,
  input  [63:0] io_out_grant_bits_data
);
  assign io_in_0_acquire_ready = io_out_acquire_ready;
  assign io_in_0_grant_valid = io_out_grant_valid;
  assign io_in_0_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_0_grant_bits_data = io_out_grant_bits_data;
  assign io_out_acquire_valid = io_in_0_acquire_valid;
  assign io_out_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign io_out_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign io_out_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign io_out_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign io_out_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign io_out_acquire_bits_union = io_in_0_acquire_bits_union;
  assign io_out_acquire_bits_data = io_in_0_acquire_bits_data;
  assign io_out_grant_ready = io_in_0_grant_ready;
endmodule
module TileLinkMemoryInterconnect(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [11:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data
);
  wire  ClientUncachedTileLinkIOArbiter_1_1_clk;
  wire  ClientUncachedTileLinkIOArbiter_1_1_reset;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_ready;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_data;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_ready;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_valid;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_data;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_ready;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_data;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_ready;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_valid;
  wire [2:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_data;
  wire [25:0] T_3009;
  ClientUncachedTileLinkIOArbiter_1 ClientUncachedTileLinkIOArbiter_1_1 (
    .clk(ClientUncachedTileLinkIOArbiter_1_1_clk),
    .reset(ClientUncachedTileLinkIOArbiter_1_1_reset),
    .io_in_0_acquire_ready(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_ready),
    .io_in_0_grant_valid(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_data),
    .io_out_acquire_ready(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_ready),
    .io_out_acquire_valid(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_valid),
    .io_out_acquire_bits_addr_block(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_block),
    .io_out_acquire_bits_client_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_client_xact_id),
    .io_out_acquire_bits_addr_beat(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_beat),
    .io_out_acquire_bits_is_builtin_type(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_is_builtin_type),
    .io_out_acquire_bits_a_type(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_a_type),
    .io_out_acquire_bits_union(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_union),
    .io_out_acquire_bits_data(ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_data),
    .io_out_grant_ready(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_ready),
    .io_out_grant_valid(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_valid),
    .io_out_grant_bits_addr_beat(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_addr_beat),
    .io_out_grant_bits_client_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_client_xact_id),
    .io_out_grant_bits_manager_xact_id(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_manager_xact_id),
    .io_out_grant_bits_is_builtin_type(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_is_builtin_type),
    .io_out_grant_bits_g_type(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_g_type),
    .io_out_grant_bits_data(ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_data)
  );
  assign io_in_0_acquire_ready = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_ready;
  assign io_in_0_grant_valid = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_valid;
  assign io_in_0_grant_bits_addr_beat = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_g_type;
  assign io_in_0_grant_bits_data = ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_bits_data;
  assign io_out_0_acquire_valid = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = T_3009;
  assign io_out_0_acquire_bits_client_xact_id = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_union;
  assign io_out_0_acquire_bits_data = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_data;
  assign io_out_0_grant_ready = ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_ready;
  assign ClientUncachedTileLinkIOArbiter_1_1_clk = clk;
  assign ClientUncachedTileLinkIOArbiter_1_1_reset = reset;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_valid = io_in_0_acquire_valid;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_union = io_in_0_acquire_bits_union;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_acquire_bits_data = io_in_0_acquire_bits_data;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_in_0_grant_ready = io_in_0_grant_ready;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_ready = io_out_0_acquire_ready;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_valid = io_out_0_grant_valid;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign ClientUncachedTileLinkIOArbiter_1_1_io_out_grant_bits_data = io_out_0_grant_bits_data;
  assign T_3009 = ClientUncachedTileLinkIOArbiter_1_1_io_out_acquire_bits_addr_block >> 1'h0;
endmodule
module LockingRRArbiter_5(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [25:0] io_in_0_bits_addr_block,
  input  [1:0] io_in_0_bits_client_xact_id,
  input  [2:0] io_in_0_bits_addr_beat,
  input   io_in_0_bits_is_builtin_type,
  input  [2:0] io_in_0_bits_a_type,
  input  [11:0] io_in_0_bits_union,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [25:0] io_in_1_bits_addr_block,
  input  [1:0] io_in_1_bits_client_xact_id,
  input  [2:0] io_in_1_bits_addr_beat,
  input   io_in_1_bits_is_builtin_type,
  input  [2:0] io_in_1_bits_a_type,
  input  [11:0] io_in_1_bits_union,
  input  [63:0] io_in_1_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [25:0] io_out_bits_addr_block,
  output [1:0] io_out_bits_client_xact_id,
  output [2:0] io_out_bits_addr_beat,
  output  io_out_bits_is_builtin_type,
  output [2:0] io_out_bits_a_type,
  output [11:0] io_out_bits_union,
  output [63:0] io_out_bits_data,
  output  io_chosen
);
  wire  choice;
  wire  GEN_0;
  wire  GEN_8;
  wire [25:0] GEN_1;
  wire [25:0] GEN_9;
  wire [1:0] GEN_2;
  wire [1:0] GEN_10;
  wire [2:0] GEN_3;
  wire [2:0] GEN_11;
  wire  GEN_4;
  wire  GEN_12;
  wire [2:0] GEN_5;
  wire [2:0] GEN_13;
  wire [11:0] GEN_6;
  wire [11:0] GEN_14;
  wire [63:0] GEN_7;
  wire [63:0] GEN_15;
  reg [2:0] T_766;
  reg [31:0] GEN_22;
  reg  T_768;
  reg [31:0] GEN_23;
  wire  T_770;
  wire [2:0] T_779_0;
  wire  T_781;
  wire  T_782;
  wire  T_783;
  wire  T_784;
  wire [3:0] T_788;
  wire [2:0] T_789;
  wire  GEN_16;
  wire [2:0] GEN_17;
  wire  GEN_18;
  reg  lastGrant;
  reg [31:0] GEN_24;
  wire  GEN_19;
  wire  T_794;
  wire  T_796;
  wire  T_799;
  wire  T_803;
  wire  T_805;
  wire  T_809;
  wire  T_811;
  wire  T_812;
  wire  T_813;
  wire  T_816;
  wire  T_817;
  wire  GEN_20;
  wire  GEN_21;
  assign io_in_0_ready = T_813;
  assign io_in_1_ready = T_817;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_block = GEN_1;
  assign io_out_bits_client_xact_id = GEN_2;
  assign io_out_bits_addr_beat = GEN_3;
  assign io_out_bits_is_builtin_type = GEN_4;
  assign io_out_bits_a_type = GEN_5;
  assign io_out_bits_union = GEN_6;
  assign io_out_bits_data = GEN_7;
  assign io_chosen = GEN_18;
  assign choice = GEN_21;
  assign GEN_0 = GEN_8;
  assign GEN_8 = io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_1 = GEN_9;
  assign GEN_9 = io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_2 = GEN_10;
  assign GEN_10 = io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_3 = GEN_11;
  assign GEN_11 = io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_4 = GEN_12;
  assign GEN_12 = io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_5 = GEN_13;
  assign GEN_13 = io_chosen ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign GEN_6 = GEN_14;
  assign GEN_14 = io_chosen ? io_in_1_bits_union : io_in_0_bits_union;
  assign GEN_7 = GEN_15;
  assign GEN_15 = io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign T_770 = T_766 != 3'h0;
  assign T_779_0 = 3'h3;
  assign T_781 = io_out_bits_a_type == T_779_0;
  assign T_782 = io_out_bits_is_builtin_type & T_781;
  assign T_783 = io_out_ready & io_out_valid;
  assign T_784 = T_783 & T_782;
  assign T_788 = T_766 + 3'h1;
  assign T_789 = T_788[2:0];
  assign GEN_16 = T_784 ? io_chosen : T_768;
  assign GEN_17 = T_784 ? T_789 : T_766;
  assign GEN_18 = T_770 ? T_768 : choice;
  assign GEN_19 = T_783 ? io_chosen : lastGrant;
  assign T_794 = 1'h1 > lastGrant;
  assign T_796 = io_in_1_valid & T_794;
  assign T_799 = T_796 | io_in_0_valid;
  assign T_803 = T_796 == 1'h0;
  assign T_805 = T_799 == 1'h0;
  assign T_809 = T_794 | T_805;
  assign T_811 = T_768 == 1'h0;
  assign T_812 = T_770 ? T_811 : T_803;
  assign T_813 = T_812 & io_out_ready;
  assign T_816 = T_770 ? T_768 : T_809;
  assign T_817 = T_816 & io_out_ready;
  assign GEN_20 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_21 = T_796 ? 1'h1 : GEN_20;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_22 = {1{$random}};
  T_766 = GEN_22[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_23 = {1{$random}};
  T_768 = GEN_23[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_24 = {1{$random}};
  lastGrant = GEN_24[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_766 <= 3'h0;
    end else begin
      if(T_784) begin
        T_766 <= T_789;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_784) begin
        T_768 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_783) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module ReorderQueue(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits_data,
  input  [1:0] io_enq_bits_tag,
  input   io_deq_valid,
  input  [1:0] io_deq_tag,
  output  io_deq_data,
  output  io_deq_matches
);
  reg  T_31 [0:3];
  reg [31:0] GEN_14;
  wire  T_31_T_47_data;
  wire [1:0] T_31_T_47_addr;
  wire  T_31_T_47_en;
  wire  T_31_T_51_data;
  wire [1:0] T_31_T_51_addr;
  wire  T_31_T_51_mask;
  wire  T_31_T_51_en;
  wire  T_41_0;
  wire  T_41_1;
  wire  T_41_2;
  wire  T_41_3;
  reg  T_45_0;
  reg [31:0] GEN_15;
  reg  T_45_1;
  reg [31:0] GEN_16;
  reg  T_45_2;
  reg [31:0] GEN_17;
  reg  T_45_3;
  reg [31:0] GEN_18;
  wire  GEN_0;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_1;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  T_49;
  wire  T_50;
  wire  GEN_2;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire  GEN_23;
  wire  GEN_3;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire  GEN_29;
  wire  GEN_30;
  wire  GEN_31;
  wire  GEN_32;
  assign io_enq_ready = GEN_0;
  assign io_deq_data = T_31_T_47_data;
  assign io_deq_matches = T_49;
  assign T_31_T_47_addr = io_deq_tag;
  assign T_31_T_47_en = 1'h1;
  assign T_31_T_47_data = T_31[T_31_T_47_addr];
  assign T_31_T_51_data = io_enq_bits_data;
  assign T_31_T_51_addr = io_enq_bits_tag;
  assign T_31_T_51_mask = T_50;
  assign T_31_T_51_en = T_50;
  assign T_41_0 = 1'h1;
  assign T_41_1 = 1'h1;
  assign T_41_2 = 1'h1;
  assign T_41_3 = 1'h1;
  assign GEN_0 = GEN_6;
  assign GEN_4 = 2'h1 == io_enq_bits_tag ? T_45_1 : T_45_0;
  assign GEN_5 = 2'h2 == io_enq_bits_tag ? T_45_2 : GEN_4;
  assign GEN_6 = 2'h3 == io_enq_bits_tag ? T_45_3 : GEN_5;
  assign GEN_1 = GEN_9;
  assign GEN_7 = 2'h1 == io_deq_tag ? T_45_1 : T_45_0;
  assign GEN_8 = 2'h2 == io_deq_tag ? T_45_2 : GEN_7;
  assign GEN_9 = 2'h3 == io_deq_tag ? T_45_3 : GEN_8;
  assign T_49 = GEN_1 == 1'h0;
  assign T_50 = io_enq_valid & io_enq_ready;
  assign GEN_2 = 1'h0;
  assign GEN_10 = 2'h0 == io_enq_bits_tag ? GEN_2 : T_45_0;
  assign GEN_11 = 2'h1 == io_enq_bits_tag ? GEN_2 : T_45_1;
  assign GEN_12 = 2'h2 == io_enq_bits_tag ? GEN_2 : T_45_2;
  assign GEN_13 = 2'h3 == io_enq_bits_tag ? GEN_2 : T_45_3;
  assign GEN_20 = T_50 ? GEN_10 : T_45_0;
  assign GEN_21 = T_50 ? GEN_11 : T_45_1;
  assign GEN_22 = T_50 ? GEN_12 : T_45_2;
  assign GEN_23 = T_50 ? GEN_13 : T_45_3;
  assign GEN_3 = 1'h1;
  assign GEN_24 = 2'h0 == io_deq_tag ? GEN_3 : GEN_20;
  assign GEN_25 = 2'h1 == io_deq_tag ? GEN_3 : GEN_21;
  assign GEN_26 = 2'h2 == io_deq_tag ? GEN_3 : GEN_22;
  assign GEN_27 = 2'h3 == io_deq_tag ? GEN_3 : GEN_23;
  assign GEN_29 = io_deq_valid ? GEN_24 : GEN_20;
  assign GEN_30 = io_deq_valid ? GEN_25 : GEN_21;
  assign GEN_31 = io_deq_valid ? GEN_26 : GEN_22;
  assign GEN_32 = io_deq_valid ? GEN_27 : GEN_23;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_14 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    T_31[initvar] = GEN_14[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_15 = {1{$random}};
  T_45_0 = GEN_15[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_16 = {1{$random}};
  T_45_1 = GEN_16[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_17 = {1{$random}};
  T_45_2 = GEN_17[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_18 = {1{$random}};
  T_45_3 = GEN_18[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(T_31_T_51_en & T_31_T_51_mask) begin
      T_31[T_31_T_51_addr] <= T_31_T_51_data;
    end
    if(reset) begin
      T_45_0 <= T_41_0;
    end else begin
      if(io_deq_valid) begin
        if(2'h0 == io_deq_tag) begin
          T_45_0 <= GEN_3;
        end else begin
          if(T_50) begin
            if(2'h0 == io_enq_bits_tag) begin
              T_45_0 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_50) begin
          if(2'h0 == io_enq_bits_tag) begin
            T_45_0 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_45_1 <= T_41_1;
    end else begin
      if(io_deq_valid) begin
        if(2'h1 == io_deq_tag) begin
          T_45_1 <= GEN_3;
        end else begin
          if(T_50) begin
            if(2'h1 == io_enq_bits_tag) begin
              T_45_1 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_50) begin
          if(2'h1 == io_enq_bits_tag) begin
            T_45_1 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_45_2 <= T_41_2;
    end else begin
      if(io_deq_valid) begin
        if(2'h2 == io_deq_tag) begin
          T_45_2 <= GEN_3;
        end else begin
          if(T_50) begin
            if(2'h2 == io_enq_bits_tag) begin
              T_45_2 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_50) begin
          if(2'h2 == io_enq_bits_tag) begin
            T_45_2 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_45_3 <= T_41_3;
    end else begin
      if(io_deq_valid) begin
        if(2'h3 == io_deq_tag) begin
          T_45_3 <= GEN_3;
        end else begin
          if(T_50) begin
            if(2'h3 == io_enq_bits_tag) begin
              T_45_3 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_50) begin
          if(2'h3 == io_enq_bits_tag) begin
            T_45_3 <= GEN_2;
          end
        end
      end
    end
  end
endmodule
module ClientTileLinkIOUnwrapper(
  input   clk,
  input   reset,
  output  io_in_acquire_ready,
  input   io_in_acquire_valid,
  input  [25:0] io_in_acquire_bits_addr_block,
  input  [1:0] io_in_acquire_bits_client_xact_id,
  input  [2:0] io_in_acquire_bits_addr_beat,
  input   io_in_acquire_bits_is_builtin_type,
  input  [2:0] io_in_acquire_bits_a_type,
  input  [11:0] io_in_acquire_bits_union,
  input  [63:0] io_in_acquire_bits_data,
  input   io_in_probe_ready,
  output  io_in_probe_valid,
  output [25:0] io_in_probe_bits_addr_block,
  output [1:0] io_in_probe_bits_p_type,
  output  io_in_release_ready,
  input   io_in_release_valid,
  input  [2:0] io_in_release_bits_addr_beat,
  input  [25:0] io_in_release_bits_addr_block,
  input  [1:0] io_in_release_bits_client_xact_id,
  input   io_in_release_bits_voluntary,
  input  [2:0] io_in_release_bits_r_type,
  input  [63:0] io_in_release_bits_data,
  input   io_in_grant_ready,
  output  io_in_grant_valid,
  output [2:0] io_in_grant_bits_addr_beat,
  output [1:0] io_in_grant_bits_client_xact_id,
  output  io_in_grant_bits_manager_xact_id,
  output  io_in_grant_bits_is_builtin_type,
  output [3:0] io_in_grant_bits_g_type,
  output [63:0] io_in_grant_bits_data,
  output  io_in_grant_bits_manager_id,
  output  io_in_finish_ready,
  input   io_in_finish_valid,
  input   io_in_finish_bits_manager_xact_id,
  input   io_in_finish_bits_manager_id,
  input   io_out_acquire_ready,
  output  io_out_acquire_valid,
  output [25:0] io_out_acquire_bits_addr_block,
  output [1:0] io_out_acquire_bits_client_xact_id,
  output [2:0] io_out_acquire_bits_addr_beat,
  output  io_out_acquire_bits_is_builtin_type,
  output [2:0] io_out_acquire_bits_a_type,
  output [11:0] io_out_acquire_bits_union,
  output [63:0] io_out_acquire_bits_data,
  output  io_out_grant_ready,
  input   io_out_grant_valid,
  input  [2:0] io_out_grant_bits_addr_beat,
  input  [1:0] io_out_grant_bits_client_xact_id,
  input   io_out_grant_bits_manager_xact_id,
  input   io_out_grant_bits_is_builtin_type,
  input  [3:0] io_out_grant_bits_g_type,
  input  [63:0] io_out_grant_bits_data
);
  wire  acqArb_clk;
  wire  acqArb_reset;
  wire  acqArb_io_in_0_ready;
  wire  acqArb_io_in_0_valid;
  wire [25:0] acqArb_io_in_0_bits_addr_block;
  wire [1:0] acqArb_io_in_0_bits_client_xact_id;
  wire [2:0] acqArb_io_in_0_bits_addr_beat;
  wire  acqArb_io_in_0_bits_is_builtin_type;
  wire [2:0] acqArb_io_in_0_bits_a_type;
  wire [11:0] acqArb_io_in_0_bits_union;
  wire [63:0] acqArb_io_in_0_bits_data;
  wire  acqArb_io_in_1_ready;
  wire  acqArb_io_in_1_valid;
  wire [25:0] acqArb_io_in_1_bits_addr_block;
  wire [1:0] acqArb_io_in_1_bits_client_xact_id;
  wire [2:0] acqArb_io_in_1_bits_addr_beat;
  wire  acqArb_io_in_1_bits_is_builtin_type;
  wire [2:0] acqArb_io_in_1_bits_a_type;
  wire [11:0] acqArb_io_in_1_bits_union;
  wire [63:0] acqArb_io_in_1_bits_data;
  wire  acqArb_io_out_ready;
  wire  acqArb_io_out_valid;
  wire [25:0] acqArb_io_out_bits_addr_block;
  wire [1:0] acqArb_io_out_bits_client_xact_id;
  wire [2:0] acqArb_io_out_bits_addr_beat;
  wire  acqArb_io_out_bits_is_builtin_type;
  wire [2:0] acqArb_io_out_bits_a_type;
  wire [11:0] acqArb_io_out_bits_union;
  wire [63:0] acqArb_io_out_bits_data;
  wire  acqArb_io_chosen;
  wire  acqRoq_clk;
  wire  acqRoq_reset;
  wire  acqRoq_io_enq_ready;
  wire  acqRoq_io_enq_valid;
  wire  acqRoq_io_enq_bits_data;
  wire [1:0] acqRoq_io_enq_bits_tag;
  wire  acqRoq_io_deq_valid;
  wire [1:0] acqRoq_io_deq_tag;
  wire  acqRoq_io_deq_data;
  wire  acqRoq_io_deq_matches;
  wire  relRoq_clk;
  wire  relRoq_reset;
  wire  relRoq_io_enq_ready;
  wire  relRoq_io_enq_valid;
  wire  relRoq_io_enq_bits_data;
  wire [1:0] relRoq_io_enq_bits_tag;
  wire  relRoq_io_deq_valid;
  wire [1:0] relRoq_io_deq_tag;
  wire  relRoq_io_deq_data;
  wire  relRoq_io_deq_matches;
  wire [2:0] T_1366_0;
  wire  T_1368;
  wire  T_1369;
  wire  T_1371;
  wire  T_1373;
  wire  acq_roq_enq;
  wire  T_1375;
  wire  T_1376;
  wire  T_1377;
  wire  T_1378;
  wire  T_1379;
  wire  T_1382;
  wire  T_1384;
  wire  rel_roq_enq;
  wire  T_1386;
  wire  acq_roq_ready;
  wire  T_1388;
  wire  rel_roq_ready;
  wire  T_1389;
  wire  T_1390;
  wire  T_1391;
  wire [2:0] T_1394;
  wire [11:0] T_1398;
  wire [25:0] T_1427_addr_block;
  wire [1:0] T_1427_client_xact_id;
  wire [2:0] T_1427_addr_beat;
  wire  T_1427_is_builtin_type;
  wire [2:0] T_1427_a_type;
  wire [11:0] T_1427_union;
  wire [63:0] T_1427_data;
  wire  T_1455;
  wire  T_1456;
  wire  T_1457;
  wire  T_1458;
  wire [25:0] T_1580_addr_block;
  wire [1:0] T_1580_client_xact_id;
  wire [2:0] T_1580_addr_beat;
  wire  T_1580_is_builtin_type;
  wire [2:0] T_1580_a_type;
  wire [11:0] T_1580_union;
  wire [63:0] T_1580_data;
  wire  T_1608;
  wire  T_1609;
  wire [2:0] T_1617_0;
  wire [3:0] GEN_0;
  wire  T_1619;
  wire  T_1620;
  wire  T_1621;
  wire  T_1624;
  wire  T_1626;
  wire  T_1627;
  wire  grant_deq_roq;
  wire  T_1628;
  wire  T_1630;
  wire  T_1631;
  wire  T_1633;
  wire  T_1634;
  wire  T_1635;
  wire  T_1636;
  wire  T_1638;
  wire [3:0] T_1639;
  wire [2:0] acq_grant_addr_beat;
  wire [1:0] acq_grant_client_xact_id;
  wire  acq_grant_manager_xact_id;
  wire  acq_grant_is_builtin_type;
  wire [3:0] acq_grant_g_type;
  wire [63:0] acq_grant_data;
  wire  T_1694;
  wire  T_1695;
  wire  T_1696;
  wire  T_1698;
  wire [2:0] rel_grant_addr_beat;
  wire [1:0] rel_grant_client_xact_id;
  wire  rel_grant_manager_xact_id;
  wire  rel_grant_is_builtin_type;
  wire [3:0] rel_grant_g_type;
  wire [63:0] rel_grant_data;
  wire [2:0] T_1754_addr_beat;
  wire [1:0] T_1754_client_xact_id;
  wire  T_1754_manager_xact_id;
  wire  T_1754_is_builtin_type;
  wire [3:0] T_1754_g_type;
  wire [63:0] T_1754_data;
  reg [25:0] GEN_1;
  reg [31:0] GEN_5;
  reg [1:0] GEN_2;
  reg [31:0] GEN_6;
  reg  GEN_3;
  reg [31:0] GEN_7;
  reg  GEN_4;
  reg [31:0] GEN_8;
  LockingRRArbiter_5 acqArb (
    .clk(acqArb_clk),
    .reset(acqArb_reset),
    .io_in_0_ready(acqArb_io_in_0_ready),
    .io_in_0_valid(acqArb_io_in_0_valid),
    .io_in_0_bits_addr_block(acqArb_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(acqArb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_addr_beat(acqArb_io_in_0_bits_addr_beat),
    .io_in_0_bits_is_builtin_type(acqArb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_a_type(acqArb_io_in_0_bits_a_type),
    .io_in_0_bits_union(acqArb_io_in_0_bits_union),
    .io_in_0_bits_data(acqArb_io_in_0_bits_data),
    .io_in_1_ready(acqArb_io_in_1_ready),
    .io_in_1_valid(acqArb_io_in_1_valid),
    .io_in_1_bits_addr_block(acqArb_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(acqArb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_addr_beat(acqArb_io_in_1_bits_addr_beat),
    .io_in_1_bits_is_builtin_type(acqArb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_a_type(acqArb_io_in_1_bits_a_type),
    .io_in_1_bits_union(acqArb_io_in_1_bits_union),
    .io_in_1_bits_data(acqArb_io_in_1_bits_data),
    .io_out_ready(acqArb_io_out_ready),
    .io_out_valid(acqArb_io_out_valid),
    .io_out_bits_addr_block(acqArb_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(acqArb_io_out_bits_client_xact_id),
    .io_out_bits_addr_beat(acqArb_io_out_bits_addr_beat),
    .io_out_bits_is_builtin_type(acqArb_io_out_bits_is_builtin_type),
    .io_out_bits_a_type(acqArb_io_out_bits_a_type),
    .io_out_bits_union(acqArb_io_out_bits_union),
    .io_out_bits_data(acqArb_io_out_bits_data),
    .io_chosen(acqArb_io_chosen)
  );
  ReorderQueue acqRoq (
    .clk(acqRoq_clk),
    .reset(acqRoq_reset),
    .io_enq_ready(acqRoq_io_enq_ready),
    .io_enq_valid(acqRoq_io_enq_valid),
    .io_enq_bits_data(acqRoq_io_enq_bits_data),
    .io_enq_bits_tag(acqRoq_io_enq_bits_tag),
    .io_deq_valid(acqRoq_io_deq_valid),
    .io_deq_tag(acqRoq_io_deq_tag),
    .io_deq_data(acqRoq_io_deq_data),
    .io_deq_matches(acqRoq_io_deq_matches)
  );
  ReorderQueue relRoq (
    .clk(relRoq_clk),
    .reset(relRoq_reset),
    .io_enq_ready(relRoq_io_enq_ready),
    .io_enq_valid(relRoq_io_enq_valid),
    .io_enq_bits_data(relRoq_io_enq_bits_data),
    .io_enq_bits_tag(relRoq_io_enq_bits_tag),
    .io_deq_valid(relRoq_io_deq_valid),
    .io_deq_tag(relRoq_io_deq_tag),
    .io_deq_data(relRoq_io_deq_data),
    .io_deq_matches(relRoq_io_deq_matches)
  );
  assign io_in_acquire_ready = T_1455;
  assign io_in_probe_valid = 1'h0;
  assign io_in_probe_bits_addr_block = GEN_1;
  assign io_in_probe_bits_p_type = GEN_2;
  assign io_in_release_ready = T_1608;
  assign io_in_grant_valid = io_out_grant_valid;
  assign io_in_grant_bits_addr_beat = T_1754_addr_beat;
  assign io_in_grant_bits_client_xact_id = T_1754_client_xact_id;
  assign io_in_grant_bits_manager_xact_id = T_1754_manager_xact_id;
  assign io_in_grant_bits_is_builtin_type = T_1754_is_builtin_type;
  assign io_in_grant_bits_g_type = T_1754_g_type;
  assign io_in_grant_bits_data = T_1754_data;
  assign io_in_grant_bits_manager_id = GEN_3;
  assign io_in_finish_ready = GEN_4;
  assign io_out_acquire_valid = acqArb_io_out_valid;
  assign io_out_acquire_bits_addr_block = acqArb_io_out_bits_addr_block;
  assign io_out_acquire_bits_client_xact_id = acqArb_io_out_bits_client_xact_id;
  assign io_out_acquire_bits_addr_beat = acqArb_io_out_bits_addr_beat;
  assign io_out_acquire_bits_is_builtin_type = acqArb_io_out_bits_is_builtin_type;
  assign io_out_acquire_bits_a_type = acqArb_io_out_bits_a_type;
  assign io_out_acquire_bits_union = acqArb_io_out_bits_union;
  assign io_out_acquire_bits_data = acqArb_io_out_bits_data;
  assign io_out_grant_ready = io_in_grant_ready;
  assign acqArb_clk = clk;
  assign acqArb_reset = reset;
  assign acqArb_io_in_0_valid = T_1391;
  assign acqArb_io_in_0_bits_addr_block = T_1427_addr_block;
  assign acqArb_io_in_0_bits_client_xact_id = T_1427_client_xact_id;
  assign acqArb_io_in_0_bits_addr_beat = T_1427_addr_beat;
  assign acqArb_io_in_0_bits_is_builtin_type = T_1427_is_builtin_type;
  assign acqArb_io_in_0_bits_a_type = T_1427_a_type;
  assign acqArb_io_in_0_bits_union = T_1427_union;
  assign acqArb_io_in_0_bits_data = T_1427_data;
  assign acqArb_io_in_1_valid = T_1458;
  assign acqArb_io_in_1_bits_addr_block = T_1580_addr_block;
  assign acqArb_io_in_1_bits_client_xact_id = T_1580_client_xact_id;
  assign acqArb_io_in_1_bits_addr_beat = T_1580_addr_beat;
  assign acqArb_io_in_1_bits_is_builtin_type = T_1580_is_builtin_type;
  assign acqArb_io_in_1_bits_a_type = T_1580_a_type;
  assign acqArb_io_in_1_bits_union = T_1580_union;
  assign acqArb_io_in_1_bits_data = T_1580_data;
  assign acqArb_io_out_ready = io_out_acquire_ready;
  assign acqRoq_clk = clk;
  assign acqRoq_reset = reset;
  assign acqRoq_io_enq_valid = T_1390;
  assign acqRoq_io_enq_bits_data = io_in_acquire_bits_is_builtin_type;
  assign acqRoq_io_enq_bits_tag = io_in_acquire_bits_client_xact_id;
  assign acqRoq_io_deq_valid = T_1628;
  assign acqRoq_io_deq_tag = io_out_grant_bits_client_xact_id;
  assign relRoq_clk = clk;
  assign relRoq_reset = reset;
  assign relRoq_io_enq_valid = T_1457;
  assign relRoq_io_enq_bits_data = io_in_release_bits_voluntary;
  assign relRoq_io_enq_bits_tag = io_in_release_bits_client_xact_id;
  assign relRoq_io_deq_valid = T_1631;
  assign relRoq_io_deq_tag = io_out_grant_bits_client_xact_id;
  assign T_1366_0 = 3'h3;
  assign T_1368 = io_in_acquire_bits_a_type == T_1366_0;
  assign T_1369 = io_in_acquire_bits_is_builtin_type & T_1368;
  assign T_1371 = T_1369 == 1'h0;
  assign T_1373 = io_in_acquire_bits_addr_beat == 3'h0;
  assign acq_roq_enq = T_1371 | T_1373;
  assign T_1375 = io_in_release_bits_r_type == 3'h0;
  assign T_1376 = io_in_release_bits_r_type == 3'h1;
  assign T_1377 = io_in_release_bits_r_type == 3'h2;
  assign T_1378 = T_1375 | T_1376;
  assign T_1379 = T_1378 | T_1377;
  assign T_1382 = T_1379 == 1'h0;
  assign T_1384 = io_in_release_bits_addr_beat == 3'h0;
  assign rel_roq_enq = T_1382 | T_1384;
  assign T_1386 = acq_roq_enq == 1'h0;
  assign acq_roq_ready = T_1386 | acqRoq_io_enq_ready;
  assign T_1388 = rel_roq_enq == 1'h0;
  assign rel_roq_ready = T_1388 | relRoq_io_enq_ready;
  assign T_1389 = io_in_acquire_valid & acqArb_io_in_0_ready;
  assign T_1390 = T_1389 & acq_roq_enq;
  assign T_1391 = io_in_acquire_valid & acq_roq_ready;
  assign T_1394 = io_in_acquire_bits_is_builtin_type ? io_in_acquire_bits_a_type : 3'h1;
  assign T_1398 = io_in_acquire_bits_is_builtin_type ? io_in_acquire_bits_union : 12'h1c1;
  assign T_1427_addr_block = io_in_acquire_bits_addr_block;
  assign T_1427_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign T_1427_addr_beat = io_in_acquire_bits_addr_beat;
  assign T_1427_is_builtin_type = 1'h1;
  assign T_1427_a_type = T_1394;
  assign T_1427_union = T_1398;
  assign T_1427_data = io_in_acquire_bits_data;
  assign T_1455 = acq_roq_ready & acqArb_io_in_0_ready;
  assign T_1456 = io_in_release_valid & acqArb_io_in_1_ready;
  assign T_1457 = T_1456 & rel_roq_enq;
  assign T_1458 = io_in_release_valid & rel_roq_ready;
  assign T_1580_addr_block = io_in_release_bits_addr_block;
  assign T_1580_client_xact_id = io_in_release_bits_client_xact_id;
  assign T_1580_addr_beat = io_in_release_bits_addr_beat;
  assign T_1580_is_builtin_type = 1'h1;
  assign T_1580_a_type = 3'h3;
  assign T_1580_union = 12'h1ff;
  assign T_1580_data = io_in_release_bits_data;
  assign T_1608 = rel_roq_ready & acqArb_io_in_1_ready;
  assign T_1609 = io_out_grant_ready & io_out_grant_valid;
  assign T_1617_0 = 3'h5;
  assign GEN_0 = {{1'd0}, T_1617_0};
  assign T_1619 = io_out_grant_bits_g_type == GEN_0;
  assign T_1620 = io_out_grant_bits_g_type == 4'h0;
  assign T_1621 = io_out_grant_bits_is_builtin_type ? T_1619 : T_1620;
  assign T_1624 = T_1621 == 1'h0;
  assign T_1626 = io_out_grant_bits_addr_beat == 3'h7;
  assign T_1627 = T_1624 | T_1626;
  assign grant_deq_roq = T_1609 & T_1627;
  assign T_1628 = acqRoq_io_deq_matches & grant_deq_roq;
  assign T_1630 = acqRoq_io_deq_matches == 1'h0;
  assign T_1631 = T_1630 & grant_deq_roq;
  assign T_1633 = grant_deq_roq == 1'h0;
  assign T_1634 = T_1633 | acqRoq_io_deq_matches;
  assign T_1635 = T_1634 | relRoq_io_deq_matches;
  assign T_1636 = T_1635 | reset;
  assign T_1638 = T_1636 == 1'h0;
  assign T_1639 = acqRoq_io_deq_data ? io_out_grant_bits_g_type : 4'h0;
  assign acq_grant_addr_beat = io_out_grant_bits_addr_beat;
  assign acq_grant_client_xact_id = io_out_grant_bits_client_xact_id;
  assign acq_grant_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign acq_grant_is_builtin_type = acqRoq_io_deq_data;
  assign acq_grant_g_type = T_1639;
  assign acq_grant_data = io_out_grant_bits_data;
  assign T_1694 = io_in_release_valid == 1'h0;
  assign T_1695 = T_1694 | io_in_release_bits_voluntary;
  assign T_1696 = T_1695 | reset;
  assign T_1698 = T_1696 == 1'h0;
  assign rel_grant_addr_beat = io_out_grant_bits_addr_beat;
  assign rel_grant_client_xact_id = io_out_grant_bits_client_xact_id;
  assign rel_grant_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign rel_grant_is_builtin_type = 1'h1;
  assign rel_grant_g_type = 4'h0;
  assign rel_grant_data = io_out_grant_bits_data;
  assign T_1754_addr_beat = acqRoq_io_deq_matches ? acq_grant_addr_beat : rel_grant_addr_beat;
  assign T_1754_client_xact_id = acqRoq_io_deq_matches ? acq_grant_client_xact_id : rel_grant_client_xact_id;
  assign T_1754_manager_xact_id = acqRoq_io_deq_matches ? acq_grant_manager_xact_id : rel_grant_manager_xact_id;
  assign T_1754_is_builtin_type = acqRoq_io_deq_matches ? acq_grant_is_builtin_type : rel_grant_is_builtin_type;
  assign T_1754_g_type = acqRoq_io_deq_matches ? acq_grant_g_type : rel_grant_g_type;
  assign T_1754_data = acqRoq_io_deq_matches ? acq_grant_data : rel_grant_data;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_5 = {1{$random}};
  GEN_1 = GEN_5[25:0];
  `endif
  `ifdef RANDOMIZE
  GEN_6 = {1{$random}};
  GEN_2 = GEN_6[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_7 = {1{$random}};
  GEN_3 = GEN_7[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_8 = {1{$random}};
  GEN_4 = GEN_8[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1638) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink Unwrapper: client_xact_id mismatch\n    at Tilelink.scala:120 assert(!grant_deq_roq || acqRoq.io.deq.matches || relRoq.io.deq.matches,\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1638) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1698) begin
          $fwrite(32'h80000002,"Assertion failed: Unwrapper can only process voluntary releases.\n    at Tilelink.scala:134 assert(!io.in.release.valid || io.in.release.bits.isVoluntary(), ---Unwrapper can only process voluntary releases.---)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1698) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module ClientTileLinkEnqueuer(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [11:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output  io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_manager_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input   io_inner_finish_bits_manager_xact_id,
  input   io_inner_finish_bits_manager_id,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [1:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [11:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [1:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [1:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id
);
  assign io_inner_acquire_ready = io_outer_acquire_ready;
  assign io_inner_probe_valid = io_outer_probe_valid;
  assign io_inner_probe_bits_addr_block = io_outer_probe_bits_addr_block;
  assign io_inner_probe_bits_p_type = io_outer_probe_bits_p_type;
  assign io_inner_release_ready = io_outer_release_ready;
  assign io_inner_grant_valid = io_outer_grant_valid;
  assign io_inner_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign io_inner_grant_bits_client_xact_id = io_outer_grant_bits_client_xact_id;
  assign io_inner_grant_bits_manager_xact_id = io_outer_grant_bits_manager_xact_id;
  assign io_inner_grant_bits_is_builtin_type = io_outer_grant_bits_is_builtin_type;
  assign io_inner_grant_bits_g_type = io_outer_grant_bits_g_type;
  assign io_inner_grant_bits_data = io_outer_grant_bits_data;
  assign io_inner_grant_bits_manager_id = io_outer_grant_bits_manager_id;
  assign io_inner_finish_ready = io_outer_finish_ready;
  assign io_outer_acquire_valid = io_inner_acquire_valid;
  assign io_outer_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign io_outer_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign io_outer_acquire_bits_union = io_inner_acquire_bits_union;
  assign io_outer_acquire_bits_data = io_inner_acquire_bits_data;
  assign io_outer_probe_ready = io_inner_probe_ready;
  assign io_outer_release_valid = io_inner_release_valid;
  assign io_outer_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign io_outer_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign io_outer_release_bits_r_type = io_inner_release_bits_r_type;
  assign io_outer_release_bits_data = io_inner_release_bits_data;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_finish_valid = io_inner_finish_valid;
  assign io_outer_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign io_outer_finish_bits_manager_id = io_inner_finish_bits_manager_id;
endmodule
module ReorderQueue_2(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [2:0] io_enq_bits_data_addr_beat,
  input   io_enq_bits_data_subblock,
  input  [1:0] io_enq_bits_tag,
  input   io_deq_valid,
  input  [1:0] io_deq_tag,
  output [2:0] io_deq_data_addr_beat,
  output  io_deq_data_subblock,
  output  io_deq_matches
);
  reg [2:0] T_229_addr_beat [0:3];
  reg [31:0] GEN_14;
  wire [2:0] T_229_addr_beat_T_245_data;
  wire [1:0] T_229_addr_beat_T_245_addr;
  wire  T_229_addr_beat_T_245_en;
  wire [2:0] T_229_addr_beat_T_271_data;
  wire [1:0] T_229_addr_beat_T_271_addr;
  wire  T_229_addr_beat_T_271_mask;
  wire  T_229_addr_beat_T_271_en;
  reg  T_229_subblock [0:3];
  reg [31:0] GEN_15;
  wire  T_229_subblock_T_245_data;
  wire [1:0] T_229_subblock_T_245_addr;
  wire  T_229_subblock_T_245_en;
  wire  T_229_subblock_T_271_data;
  wire [1:0] T_229_subblock_T_271_addr;
  wire  T_229_subblock_T_271_mask;
  wire  T_229_subblock_T_271_en;
  wire  T_239_0;
  wire  T_239_1;
  wire  T_239_2;
  wire  T_239_3;
  reg  T_243_0;
  reg [31:0] GEN_16;
  reg  T_243_1;
  reg [31:0] GEN_17;
  reg  T_243_2;
  reg [31:0] GEN_18;
  reg  T_243_3;
  reg [31:0] GEN_19;
  wire  GEN_0;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_1;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  T_269;
  wire  T_270;
  wire  GEN_2;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_3;
  wire  GEN_26;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_29;
  wire  GEN_31;
  wire  GEN_32;
  wire  GEN_33;
  wire  GEN_34;
  assign io_enq_ready = GEN_0;
  assign io_deq_data_addr_beat = T_229_addr_beat_T_245_data;
  assign io_deq_data_subblock = T_229_subblock_T_245_data;
  assign io_deq_matches = T_269;
  assign T_229_addr_beat_T_245_addr = io_deq_tag;
  assign T_229_addr_beat_T_245_en = 1'h1;
  assign T_229_addr_beat_T_245_data = T_229_addr_beat[T_229_addr_beat_T_245_addr];
  assign T_229_addr_beat_T_271_data = io_enq_bits_data_addr_beat;
  assign T_229_addr_beat_T_271_addr = io_enq_bits_tag;
  assign T_229_addr_beat_T_271_mask = T_270;
  assign T_229_addr_beat_T_271_en = T_270;
  assign T_229_subblock_T_245_addr = io_deq_tag;
  assign T_229_subblock_T_245_en = 1'h1;
  assign T_229_subblock_T_245_data = T_229_subblock[T_229_subblock_T_245_addr];
  assign T_229_subblock_T_271_data = io_enq_bits_data_subblock;
  assign T_229_subblock_T_271_addr = io_enq_bits_tag;
  assign T_229_subblock_T_271_mask = T_270;
  assign T_229_subblock_T_271_en = T_270;
  assign T_239_0 = 1'h1;
  assign T_239_1 = 1'h1;
  assign T_239_2 = 1'h1;
  assign T_239_3 = 1'h1;
  assign GEN_0 = GEN_6;
  assign GEN_4 = 2'h1 == io_enq_bits_tag ? T_243_1 : T_243_0;
  assign GEN_5 = 2'h2 == io_enq_bits_tag ? T_243_2 : GEN_4;
  assign GEN_6 = 2'h3 == io_enq_bits_tag ? T_243_3 : GEN_5;
  assign GEN_1 = GEN_9;
  assign GEN_7 = 2'h1 == io_deq_tag ? T_243_1 : T_243_0;
  assign GEN_8 = 2'h2 == io_deq_tag ? T_243_2 : GEN_7;
  assign GEN_9 = 2'h3 == io_deq_tag ? T_243_3 : GEN_8;
  assign T_269 = GEN_1 == 1'h0;
  assign T_270 = io_enq_valid & io_enq_ready;
  assign GEN_2 = 1'h0;
  assign GEN_10 = 2'h0 == io_enq_bits_tag ? GEN_2 : T_243_0;
  assign GEN_11 = 2'h1 == io_enq_bits_tag ? GEN_2 : T_243_1;
  assign GEN_12 = 2'h2 == io_enq_bits_tag ? GEN_2 : T_243_2;
  assign GEN_13 = 2'h3 == io_enq_bits_tag ? GEN_2 : T_243_3;
  assign GEN_22 = T_270 ? GEN_10 : T_243_0;
  assign GEN_23 = T_270 ? GEN_11 : T_243_1;
  assign GEN_24 = T_270 ? GEN_12 : T_243_2;
  assign GEN_25 = T_270 ? GEN_13 : T_243_3;
  assign GEN_3 = 1'h1;
  assign GEN_26 = 2'h0 == io_deq_tag ? GEN_3 : GEN_22;
  assign GEN_27 = 2'h1 == io_deq_tag ? GEN_3 : GEN_23;
  assign GEN_28 = 2'h2 == io_deq_tag ? GEN_3 : GEN_24;
  assign GEN_29 = 2'h3 == io_deq_tag ? GEN_3 : GEN_25;
  assign GEN_31 = io_deq_valid ? GEN_26 : GEN_22;
  assign GEN_32 = io_deq_valid ? GEN_27 : GEN_23;
  assign GEN_33 = io_deq_valid ? GEN_28 : GEN_24;
  assign GEN_34 = io_deq_valid ? GEN_29 : GEN_25;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_14 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    T_229_addr_beat[initvar] = GEN_14[2:0];
  `endif
  GEN_15 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    T_229_subblock[initvar] = GEN_15[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_16 = {1{$random}};
  T_243_0 = GEN_16[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_17 = {1{$random}};
  T_243_1 = GEN_17[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_18 = {1{$random}};
  T_243_2 = GEN_18[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_19 = {1{$random}};
  T_243_3 = GEN_19[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(T_229_addr_beat_T_271_en & T_229_addr_beat_T_271_mask) begin
      T_229_addr_beat[T_229_addr_beat_T_271_addr] <= T_229_addr_beat_T_271_data;
    end
    if(T_229_subblock_T_271_en & T_229_subblock_T_271_mask) begin
      T_229_subblock[T_229_subblock_T_271_addr] <= T_229_subblock_T_271_data;
    end
    if(reset) begin
      T_243_0 <= T_239_0;
    end else begin
      if(io_deq_valid) begin
        if(2'h0 == io_deq_tag) begin
          T_243_0 <= GEN_3;
        end else begin
          if(T_270) begin
            if(2'h0 == io_enq_bits_tag) begin
              T_243_0 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_270) begin
          if(2'h0 == io_enq_bits_tag) begin
            T_243_0 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_243_1 <= T_239_1;
    end else begin
      if(io_deq_valid) begin
        if(2'h1 == io_deq_tag) begin
          T_243_1 <= GEN_3;
        end else begin
          if(T_270) begin
            if(2'h1 == io_enq_bits_tag) begin
              T_243_1 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_270) begin
          if(2'h1 == io_enq_bits_tag) begin
            T_243_1 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_243_2 <= T_239_2;
    end else begin
      if(io_deq_valid) begin
        if(2'h2 == io_deq_tag) begin
          T_243_2 <= GEN_3;
        end else begin
          if(T_270) begin
            if(2'h2 == io_enq_bits_tag) begin
              T_243_2 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_270) begin
          if(2'h2 == io_enq_bits_tag) begin
            T_243_2 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_243_3 <= T_239_3;
    end else begin
      if(io_deq_valid) begin
        if(2'h3 == io_deq_tag) begin
          T_243_3 <= GEN_3;
        end else begin
          if(T_270) begin
            if(2'h3 == io_enq_bits_tag) begin
              T_243_3 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_270) begin
          if(2'h3 == io_enq_bits_tag) begin
            T_243_3 <= GEN_2;
          end
        end
      end
    end
  end
endmodule
module IdMapper(
  input   clk,
  input   reset,
  input   io_req_valid,
  output  io_req_ready,
  input  [1:0] io_req_in_id,
  output [4:0] io_req_out_id,
  input   io_resp_valid,
  output  io_resp_matches,
  input  [4:0] io_resp_out_id,
  output [1:0] io_resp_in_id
);
  assign io_req_ready = 1'h1;
  assign io_req_out_id = {{3'd0}, io_req_in_id};
  assign io_resp_matches = 1'h1;
  assign io_resp_in_id = io_resp_out_id[1:0];
endmodule
module LockingArbiter(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  input   io_in_0_bits_client_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [1:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_is_builtin_type,
  input  [3:0] io_in_1_bits_g_type,
  input  [63:0] io_in_1_bits_data,
  input   io_in_1_bits_client_id,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_out_bits_client_id,
  output  io_chosen
);
  wire  choice;
  wire  GEN_0;
  wire  GEN_8;
  wire [2:0] GEN_1;
  wire [2:0] GEN_9;
  wire [1:0] GEN_2;
  wire [1:0] GEN_10;
  wire  GEN_3;
  wire  GEN_11;
  wire  GEN_4;
  wire  GEN_12;
  wire [3:0] GEN_5;
  wire [3:0] GEN_13;
  wire [63:0] GEN_6;
  wire [63:0] GEN_14;
  wire  GEN_7;
  wire  GEN_15;
  reg [2:0] T_766;
  reg [31:0] GEN_21;
  reg  T_768;
  reg [31:0] GEN_22;
  wire  T_770;
  wire [2:0] T_778_0;
  wire [3:0] GEN_20;
  wire  T_780;
  wire  T_781;
  wire  T_782;
  wire  T_784;
  wire  T_785;
  wire [3:0] T_789;
  wire [2:0] T_790;
  wire  GEN_16;
  wire [2:0] GEN_17;
  wire  GEN_18;
  wire  T_793;
  wire  T_795;
  wire  T_796;
  wire  T_797;
  wire  T_800;
  wire  T_801;
  wire  GEN_19;
  assign io_in_0_ready = T_797;
  assign io_in_1_ready = T_801;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_beat = GEN_1;
  assign io_out_bits_client_xact_id = GEN_2;
  assign io_out_bits_manager_xact_id = GEN_3;
  assign io_out_bits_is_builtin_type = GEN_4;
  assign io_out_bits_g_type = GEN_5;
  assign io_out_bits_data = GEN_6;
  assign io_out_bits_client_id = GEN_7;
  assign io_chosen = GEN_18;
  assign choice = GEN_19;
  assign GEN_0 = GEN_8;
  assign GEN_8 = io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_1 = GEN_9;
  assign GEN_9 = io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_2 = GEN_10;
  assign GEN_10 = io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_3 = GEN_11;
  assign GEN_11 = io_chosen ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign GEN_4 = GEN_12;
  assign GEN_12 = io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_5 = GEN_13;
  assign GEN_13 = io_chosen ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign GEN_6 = GEN_14;
  assign GEN_14 = io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_7 = GEN_15;
  assign GEN_15 = io_chosen ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign T_770 = T_766 != 3'h0;
  assign T_778_0 = 3'h5;
  assign GEN_20 = {{1'd0}, T_778_0};
  assign T_780 = io_out_bits_g_type == GEN_20;
  assign T_781 = io_out_bits_g_type == 4'h0;
  assign T_782 = io_out_bits_is_builtin_type ? T_780 : T_781;
  assign T_784 = io_out_ready & io_out_valid;
  assign T_785 = T_784 & T_782;
  assign T_789 = T_766 + 3'h1;
  assign T_790 = T_789[2:0];
  assign GEN_16 = T_785 ? io_chosen : T_768;
  assign GEN_17 = T_785 ? T_790 : T_766;
  assign GEN_18 = T_770 ? T_768 : choice;
  assign T_793 = io_in_0_valid == 1'h0;
  assign T_795 = T_768 == 1'h0;
  assign T_796 = T_770 ? T_795 : 1'h1;
  assign T_797 = T_796 & io_out_ready;
  assign T_800 = T_770 ? T_768 : T_793;
  assign T_801 = T_800 & io_out_ready;
  assign GEN_19 = io_in_0_valid ? 1'h0 : 1'h1;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_21 = {1{$random}};
  T_766 = GEN_21[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_22 = {1{$random}};
  T_768 = GEN_22[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_766 <= 3'h0;
    end else begin
      if(T_785) begin
        T_766 <= T_790;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_785) begin
        T_768 <= io_chosen;
      end
    end
  end
endmodule
module NastiIOTileLinkIOConverter(
  input   clk,
  input   reset,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [11:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data,
  input   io_nasti_aw_ready,
  output  io_nasti_aw_valid,
  output [31:0] io_nasti_aw_bits_addr,
  output [7:0] io_nasti_aw_bits_len,
  output [2:0] io_nasti_aw_bits_size,
  output [1:0] io_nasti_aw_bits_burst,
  output  io_nasti_aw_bits_lock,
  output [3:0] io_nasti_aw_bits_cache,
  output [2:0] io_nasti_aw_bits_prot,
  output [3:0] io_nasti_aw_bits_qos,
  output [3:0] io_nasti_aw_bits_region,
  output [4:0] io_nasti_aw_bits_id,
  output  io_nasti_aw_bits_user,
  input   io_nasti_w_ready,
  output  io_nasti_w_valid,
  output [63:0] io_nasti_w_bits_data,
  output  io_nasti_w_bits_last,
  output [4:0] io_nasti_w_bits_id,
  output [7:0] io_nasti_w_bits_strb,
  output  io_nasti_w_bits_user,
  output  io_nasti_b_ready,
  input   io_nasti_b_valid,
  input  [1:0] io_nasti_b_bits_resp,
  input  [4:0] io_nasti_b_bits_id,
  input   io_nasti_b_bits_user,
  input   io_nasti_ar_ready,
  output  io_nasti_ar_valid,
  output [31:0] io_nasti_ar_bits_addr,
  output [7:0] io_nasti_ar_bits_len,
  output [2:0] io_nasti_ar_bits_size,
  output [1:0] io_nasti_ar_bits_burst,
  output  io_nasti_ar_bits_lock,
  output [3:0] io_nasti_ar_bits_cache,
  output [2:0] io_nasti_ar_bits_prot,
  output [3:0] io_nasti_ar_bits_qos,
  output [3:0] io_nasti_ar_bits_region,
  output [4:0] io_nasti_ar_bits_id,
  output  io_nasti_ar_bits_user,
  output  io_nasti_r_ready,
  input   io_nasti_r_valid,
  input  [1:0] io_nasti_r_bits_resp,
  input  [63:0] io_nasti_r_bits_data,
  input   io_nasti_r_bits_last,
  input  [4:0] io_nasti_r_bits_id,
  input   io_nasti_r_bits_user
);
  wire [2:0] T_688_0;
  wire [2:0] T_688_1;
  wire [2:0] T_688_2;
  wire  T_690;
  wire  T_691;
  wire  T_692;
  wire  T_693;
  wire  T_694;
  wire  has_data;
  wire [2:0] T_703_0;
  wire [2:0] T_703_1;
  wire [2:0] T_703_2;
  wire  T_705;
  wire  T_706;
  wire  T_707;
  wire  T_708;
  wire  T_709;
  wire  is_subblock;
  wire [2:0] T_718_0;
  wire  T_720;
  wire  is_multibeat;
  wire  T_721;
  wire  T_722;
  reg [2:0] tl_cnt_out;
  reg [31:0] GEN_11;
  wire  T_725;
  wire [3:0] T_727;
  wire [2:0] T_728;
  wire [2:0] GEN_0;
  wire  tl_wrap_out;
  wire  T_730;
  wire  get_valid;
  wire  put_valid;
  wire  roq_clk;
  wire  roq_reset;
  wire  roq_io_enq_ready;
  wire  roq_io_enq_valid;
  wire [2:0] roq_io_enq_bits_data_addr_beat;
  wire  roq_io_enq_bits_data_subblock;
  wire [1:0] roq_io_enq_bits_tag;
  wire  roq_io_deq_valid;
  wire [1:0] roq_io_deq_tag;
  wire [2:0] roq_io_deq_data_addr_beat;
  wire  roq_io_deq_data_subblock;
  wire  roq_io_deq_matches;
  wire  get_id_mapper_clk;
  wire  get_id_mapper_reset;
  wire  get_id_mapper_io_req_valid;
  wire  get_id_mapper_io_req_ready;
  wire [1:0] get_id_mapper_io_req_in_id;
  wire [4:0] get_id_mapper_io_req_out_id;
  wire  get_id_mapper_io_resp_valid;
  wire  get_id_mapper_io_resp_matches;
  wire [4:0] get_id_mapper_io_resp_out_id;
  wire [1:0] get_id_mapper_io_resp_in_id;
  wire  put_id_mapper_clk;
  wire  put_id_mapper_reset;
  wire  put_id_mapper_io_req_valid;
  wire  put_id_mapper_io_req_ready;
  wire [1:0] put_id_mapper_io_req_in_id;
  wire [4:0] put_id_mapper_io_req_out_id;
  wire  put_id_mapper_io_resp_valid;
  wire  put_id_mapper_io_resp_matches;
  wire [4:0] put_id_mapper_io_resp_out_id;
  wire [1:0] put_id_mapper_io_resp_in_id;
  wire  T_755;
  wire  put_id_mask;
  wire  T_757;
  wire  put_id_ready;
  reg  w_inflight;
  reg [31:0] GEN_12;
  reg [4:0] w_id;
  reg [31:0] GEN_13;
  wire  aw_ready;
  wire  T_760;
  wire  T_762;
  wire  T_763;
  reg [2:0] nasti_cnt_out;
  reg [31:0] GEN_14;
  wire  T_766;
  wire [3:0] T_768;
  wire [2:0] T_769;
  wire [2:0] GEN_1;
  wire  nasti_wrap_out;
  wire  T_770;
  wire  T_771;
  wire  T_773;
  wire  T_774;
  wire  T_775;
  wire  T_776;
  wire  T_778;
  wire  T_779;
  wire  T_780;
  wire  T_781;
  wire  T_782;
  wire  T_784;
  wire [2:0] T_792_0;
  wire [2:0] T_792_1;
  wire  T_794;
  wire  T_795;
  wire  T_796;
  wire  T_797;
  wire [2:0] T_798;
  wire [2:0] T_800;
  wire [28:0] T_801;
  wire [31:0] T_802;
  wire [2:0] T_803;
  wire  T_813;
  wire [2:0] T_814;
  wire  T_815;
  wire [2:0] T_816;
  wire  T_817;
  wire [2:0] T_818;
  wire  T_819;
  wire [2:0] T_820;
  wire  T_821;
  wire [2:0] T_822;
  wire  T_823;
  wire [2:0] T_824;
  wire  T_825;
  wire [2:0] T_826;
  wire  T_827;
  wire [2:0] T_828;
  wire [2:0] T_830;
  wire [2:0] T_833;
  wire [31:0] T_853_addr;
  wire [7:0] T_853_len;
  wire [2:0] T_853_size;
  wire [1:0] T_853_burst;
  wire  T_853_lock;
  wire [3:0] T_853_cache;
  wire [2:0] T_853_prot;
  wire [3:0] T_853_qos;
  wire [3:0] T_853_region;
  wire [4:0] T_853_id;
  wire  T_853_user;
  wire  T_872;
  wire  T_873;
  wire  T_875;
  wire [1:0] T_877;
  wire  T_878;
  wire  T_879;
  wire [3:0] T_883;
  wire [3:0] T_887;
  wire [7:0] T_888;
  wire  T_890;
  wire  T_891;
  wire  T_893;
  wire  T_894;
  wire  T_895;
  wire [7:0] T_896;
  wire [7:0] T_898;
  wire [7:0] T_899;
  wire [7:0] T_900;
  wire  T_901;
  wire  T_902;
  wire  T_903;
  wire  T_904;
  wire  T_905;
  wire  T_906;
  wire  T_907;
  wire  T_908;
  wire  T_909;
  wire  T_910;
  wire  T_911;
  wire  T_912;
  wire  T_913;
  wire  T_914;
  wire  T_921;
  wire [1:0] T_922;
  wire [1:0] T_924;
  wire  T_925;
  wire  T_926;
  wire  T_927;
  wire  T_928;
  wire  T_929;
  wire  T_930;
  wire  T_931;
  wire  T_932;
  wire [2:0] T_933;
  wire [1:0] T_935;
  wire  T_936;
  wire  T_937;
  wire  T_938;
  wire  T_939;
  wire  T_940;
  wire  T_941;
  wire  T_942;
  wire  T_943;
  wire  T_944;
  wire  T_945;
  wire  T_946;
  wire  T_947;
  wire  T_948;
  wire  T_949;
  wire  T_950;
  wire  T_951;
  wire  T_952;
  wire  T_953;
  wire [3:0] put_offset;
  wire [1:0] put_size;
  wire  T_956;
  wire  T_957;
  wire  T_958;
  wire  T_959;
  wire [2:0] T_967_0;
  wire [2:0] T_967_1;
  wire  T_969;
  wire  T_970;
  wire  T_971;
  wire  T_972;
  wire [2:0] T_975;
  wire [31:0] T_977;
  wire [3:0] T_979;
  wire [31:0] GEN_7;
  wire [31:0] T_980;
  wire [1:0] T_982;
  wire [2:0] T_985;
  wire [31:0] T_998_addr;
  wire [7:0] T_998_len;
  wire [2:0] T_998_size;
  wire [1:0] T_998_burst;
  wire  T_998_lock;
  wire [3:0] T_998_cache;
  wire [2:0] T_998_prot;
  wire [3:0] T_998_qos;
  wire [3:0] T_998_region;
  wire [4:0] T_998_id;
  wire  T_998_user;
  wire  T_1017;
  wire  T_1050;
  wire  T_1051;
  wire [63:0] T_1058_data;
  wire  T_1058_last;
  wire [4:0] T_1058_id;
  wire [7:0] T_1058_strb;
  wire  T_1058_user;
  wire  T_1065;
  wire  T_1066;
  wire  T_1067;
  wire  T_1068;
  wire  T_1069;
  wire  T_1073;
  wire  T_1074;
  wire  GEN_2;
  wire [4:0] GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire  T_1077;
  wire [2:0] T_1085_0;
  wire [3:0] GEN_8;
  wire  T_1087;
  wire  T_1088;
  wire  T_1089;
  wire  T_1091;
  reg [2:0] tl_cnt_in;
  reg [31:0] GEN_15;
  wire [3:0] T_1096;
  wire [2:0] T_1097;
  wire [2:0] GEN_6;
  wire  gnt_arb_clk;
  wire  gnt_arb_reset;
  wire  gnt_arb_io_in_0_ready;
  wire  gnt_arb_io_in_0_valid;
  wire [2:0] gnt_arb_io_in_0_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_0_bits_client_xact_id;
  wire  gnt_arb_io_in_0_bits_manager_xact_id;
  wire  gnt_arb_io_in_0_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_0_bits_g_type;
  wire [63:0] gnt_arb_io_in_0_bits_data;
  wire  gnt_arb_io_in_0_bits_client_id;
  wire  gnt_arb_io_in_1_ready;
  wire  gnt_arb_io_in_1_valid;
  wire [2:0] gnt_arb_io_in_1_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_1_bits_client_xact_id;
  wire  gnt_arb_io_in_1_bits_manager_xact_id;
  wire  gnt_arb_io_in_1_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_1_bits_g_type;
  wire [63:0] gnt_arb_io_in_1_bits_data;
  wire  gnt_arb_io_in_1_bits_client_id;
  wire  gnt_arb_io_out_ready;
  wire  gnt_arb_io_out_valid;
  wire [2:0] gnt_arb_io_out_bits_addr_beat;
  wire [1:0] gnt_arb_io_out_bits_client_xact_id;
  wire  gnt_arb_io_out_bits_manager_xact_id;
  wire  gnt_arb_io_out_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_out_bits_g_type;
  wire [63:0] gnt_arb_io_out_bits_data;
  wire  gnt_arb_io_out_bits_client_id;
  wire  gnt_arb_io_chosen;
  wire [2:0] T_1129;
  wire [2:0] T_1131;
  wire [2:0] T_1159_addr_beat;
  wire [1:0] T_1159_client_xact_id;
  wire  T_1159_manager_xact_id;
  wire  T_1159_is_builtin_type;
  wire [3:0] T_1159_g_type;
  wire [63:0] T_1159_data;
  wire  T_1187;
  wire  T_1188;
  wire  T_1189;
  wire  T_1191;
  wire  T_1193;
  wire  T_1194;
  wire  T_1195;
  wire  T_1197;
  wire [2:0] T_1230_addr_beat;
  wire [1:0] T_1230_client_xact_id;
  wire  T_1230_manager_xact_id;
  wire  T_1230_is_builtin_type;
  wire [3:0] T_1230_g_type;
  wire [63:0] T_1230_data;
  wire  T_1258;
  wire  T_1259;
  wire  T_1260;
  wire  T_1262;
  wire  T_1264;
  wire  T_1266;
  wire  T_1267;
  wire  T_1268;
  wire  T_1270;
  wire  T_1272;
  wire  T_1274;
  wire  T_1275;
  wire  T_1276;
  wire  T_1278;
  reg  GEN_9;
  reg [31:0] GEN_16;
  reg  GEN_10;
  reg [31:0] GEN_17;
  ReorderQueue_2 roq (
    .clk(roq_clk),
    .reset(roq_reset),
    .io_enq_ready(roq_io_enq_ready),
    .io_enq_valid(roq_io_enq_valid),
    .io_enq_bits_data_addr_beat(roq_io_enq_bits_data_addr_beat),
    .io_enq_bits_data_subblock(roq_io_enq_bits_data_subblock),
    .io_enq_bits_tag(roq_io_enq_bits_tag),
    .io_deq_valid(roq_io_deq_valid),
    .io_deq_tag(roq_io_deq_tag),
    .io_deq_data_addr_beat(roq_io_deq_data_addr_beat),
    .io_deq_data_subblock(roq_io_deq_data_subblock),
    .io_deq_matches(roq_io_deq_matches)
  );
  IdMapper get_id_mapper (
    .clk(get_id_mapper_clk),
    .reset(get_id_mapper_reset),
    .io_req_valid(get_id_mapper_io_req_valid),
    .io_req_ready(get_id_mapper_io_req_ready),
    .io_req_in_id(get_id_mapper_io_req_in_id),
    .io_req_out_id(get_id_mapper_io_req_out_id),
    .io_resp_valid(get_id_mapper_io_resp_valid),
    .io_resp_matches(get_id_mapper_io_resp_matches),
    .io_resp_out_id(get_id_mapper_io_resp_out_id),
    .io_resp_in_id(get_id_mapper_io_resp_in_id)
  );
  IdMapper put_id_mapper (
    .clk(put_id_mapper_clk),
    .reset(put_id_mapper_reset),
    .io_req_valid(put_id_mapper_io_req_valid),
    .io_req_ready(put_id_mapper_io_req_ready),
    .io_req_in_id(put_id_mapper_io_req_in_id),
    .io_req_out_id(put_id_mapper_io_req_out_id),
    .io_resp_valid(put_id_mapper_io_resp_valid),
    .io_resp_matches(put_id_mapper_io_resp_matches),
    .io_resp_out_id(put_id_mapper_io_resp_out_id),
    .io_resp_in_id(put_id_mapper_io_resp_in_id)
  );
  LockingArbiter gnt_arb (
    .clk(gnt_arb_clk),
    .reset(gnt_arb_reset),
    .io_in_0_ready(gnt_arb_io_in_0_ready),
    .io_in_0_valid(gnt_arb_io_in_0_valid),
    .io_in_0_bits_addr_beat(gnt_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(gnt_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(gnt_arb_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(gnt_arb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(gnt_arb_io_in_0_bits_g_type),
    .io_in_0_bits_data(gnt_arb_io_in_0_bits_data),
    .io_in_0_bits_client_id(gnt_arb_io_in_0_bits_client_id),
    .io_in_1_ready(gnt_arb_io_in_1_ready),
    .io_in_1_valid(gnt_arb_io_in_1_valid),
    .io_in_1_bits_addr_beat(gnt_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_client_xact_id(gnt_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_manager_xact_id(gnt_arb_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_is_builtin_type(gnt_arb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_g_type(gnt_arb_io_in_1_bits_g_type),
    .io_in_1_bits_data(gnt_arb_io_in_1_bits_data),
    .io_in_1_bits_client_id(gnt_arb_io_in_1_bits_client_id),
    .io_out_ready(gnt_arb_io_out_ready),
    .io_out_valid(gnt_arb_io_out_valid),
    .io_out_bits_addr_beat(gnt_arb_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(gnt_arb_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(gnt_arb_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(gnt_arb_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(gnt_arb_io_out_bits_g_type),
    .io_out_bits_data(gnt_arb_io_out_bits_data),
    .io_out_bits_client_id(gnt_arb_io_out_bits_client_id),
    .io_chosen(gnt_arb_io_chosen)
  );
  assign io_tl_acquire_ready = T_1069;
  assign io_tl_grant_valid = gnt_arb_io_out_valid;
  assign io_tl_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_tl_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_tl_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_tl_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_nasti_aw_valid = T_959;
  assign io_nasti_aw_bits_addr = T_998_addr;
  assign io_nasti_aw_bits_len = T_998_len;
  assign io_nasti_aw_bits_size = T_998_size;
  assign io_nasti_aw_bits_burst = T_998_burst;
  assign io_nasti_aw_bits_lock = T_998_lock;
  assign io_nasti_aw_bits_cache = T_998_cache;
  assign io_nasti_aw_bits_prot = T_998_prot;
  assign io_nasti_aw_bits_qos = T_998_qos;
  assign io_nasti_aw_bits_region = T_998_region;
  assign io_nasti_aw_bits_id = T_998_id;
  assign io_nasti_aw_bits_user = T_998_user;
  assign io_nasti_w_valid = T_1017;
  assign io_nasti_w_bits_data = T_1058_data;
  assign io_nasti_w_bits_last = T_1058_last;
  assign io_nasti_w_bits_id = T_1058_id;
  assign io_nasti_w_bits_strb = T_1058_strb;
  assign io_nasti_w_bits_user = T_1058_user;
  assign io_nasti_b_ready = gnt_arb_io_in_1_ready;
  assign io_nasti_ar_valid = T_784;
  assign io_nasti_ar_bits_addr = T_853_addr;
  assign io_nasti_ar_bits_len = T_853_len;
  assign io_nasti_ar_bits_size = T_853_size;
  assign io_nasti_ar_bits_burst = T_853_burst;
  assign io_nasti_ar_bits_lock = T_853_lock;
  assign io_nasti_ar_bits_cache = T_853_cache;
  assign io_nasti_ar_bits_prot = T_853_prot;
  assign io_nasti_ar_bits_qos = T_853_qos;
  assign io_nasti_ar_bits_region = T_853_region;
  assign io_nasti_ar_bits_id = T_853_id;
  assign io_nasti_ar_bits_user = T_853_user;
  assign io_nasti_r_ready = gnt_arb_io_in_0_ready;
  assign T_688_0 = 3'h2;
  assign T_688_1 = 3'h3;
  assign T_688_2 = 3'h4;
  assign T_690 = io_tl_acquire_bits_a_type == T_688_0;
  assign T_691 = io_tl_acquire_bits_a_type == T_688_1;
  assign T_692 = io_tl_acquire_bits_a_type == T_688_2;
  assign T_693 = T_690 | T_691;
  assign T_694 = T_693 | T_692;
  assign has_data = io_tl_acquire_bits_is_builtin_type & T_694;
  assign T_703_0 = 3'h2;
  assign T_703_1 = 3'h0;
  assign T_703_2 = 3'h4;
  assign T_705 = io_tl_acquire_bits_a_type == T_703_0;
  assign T_706 = io_tl_acquire_bits_a_type == T_703_1;
  assign T_707 = io_tl_acquire_bits_a_type == T_703_2;
  assign T_708 = T_705 | T_706;
  assign T_709 = T_708 | T_707;
  assign is_subblock = io_tl_acquire_bits_is_builtin_type & T_709;
  assign T_718_0 = 3'h3;
  assign T_720 = io_tl_acquire_bits_a_type == T_718_0;
  assign is_multibeat = io_tl_acquire_bits_is_builtin_type & T_720;
  assign T_721 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign T_722 = T_721 & is_multibeat;
  assign T_725 = tl_cnt_out == 3'h7;
  assign T_727 = tl_cnt_out + 3'h1;
  assign T_728 = T_727[2:0];
  assign GEN_0 = T_722 ? T_728 : tl_cnt_out;
  assign tl_wrap_out = T_722 & T_725;
  assign T_730 = has_data == 1'h0;
  assign get_valid = io_tl_acquire_valid & T_730;
  assign put_valid = io_tl_acquire_valid & has_data;
  assign roq_clk = clk;
  assign roq_reset = reset;
  assign roq_io_enq_valid = T_771;
  assign roq_io_enq_bits_data_addr_beat = io_tl_acquire_bits_addr_beat;
  assign roq_io_enq_bits_data_subblock = is_subblock;
  assign roq_io_enq_bits_tag = io_nasti_ar_bits_id[1:0];
  assign roq_io_deq_valid = T_774;
  assign roq_io_deq_tag = io_nasti_r_bits_id[1:0];
  assign get_id_mapper_clk = clk;
  assign get_id_mapper_reset = reset;
  assign get_id_mapper_io_req_valid = T_776;
  assign get_id_mapper_io_req_in_id = io_tl_acquire_bits_client_xact_id;
  assign get_id_mapper_io_resp_valid = T_778;
  assign get_id_mapper_io_resp_out_id = io_nasti_r_bits_id;
  assign put_id_mapper_clk = clk;
  assign put_id_mapper_reset = reset;
  assign put_id_mapper_io_req_valid = T_781;
  assign put_id_mapper_io_req_in_id = io_tl_acquire_bits_client_xact_id;
  assign put_id_mapper_io_resp_valid = T_782;
  assign put_id_mapper_io_resp_out_id = io_nasti_b_bits_id;
  assign T_755 = io_tl_acquire_bits_addr_beat == 3'h0;
  assign put_id_mask = is_subblock | T_755;
  assign T_757 = put_id_mask == 1'h0;
  assign put_id_ready = put_id_mapper_io_req_ready | T_757;
  assign aw_ready = w_inflight | io_nasti_aw_ready;
  assign T_760 = io_nasti_r_ready & io_nasti_r_valid;
  assign T_762 = roq_io_deq_data_subblock == 1'h0;
  assign T_763 = T_760 & T_762;
  assign T_766 = nasti_cnt_out == 3'h7;
  assign T_768 = nasti_cnt_out + 3'h1;
  assign T_769 = T_768[2:0];
  assign GEN_1 = T_763 ? T_769 : nasti_cnt_out;
  assign nasti_wrap_out = T_763 & T_766;
  assign T_770 = get_valid & io_nasti_ar_ready;
  assign T_771 = T_770 & get_id_mapper_io_req_ready;
  assign T_773 = nasti_wrap_out | roq_io_deq_data_subblock;
  assign T_774 = T_760 & T_773;
  assign T_775 = get_valid & roq_io_enq_ready;
  assign T_776 = T_775 & io_nasti_ar_ready;
  assign T_778 = T_760 & io_nasti_r_bits_last;
  assign T_779 = put_valid & aw_ready;
  assign T_780 = T_779 & io_nasti_w_ready;
  assign T_781 = T_780 & put_id_mask;
  assign T_782 = io_nasti_b_ready & io_nasti_b_valid;
  assign T_784 = T_775 & get_id_mapper_io_req_ready;
  assign T_792_0 = 3'h0;
  assign T_792_1 = 3'h4;
  assign T_794 = io_tl_acquire_bits_a_type == T_792_0;
  assign T_795 = io_tl_acquire_bits_a_type == T_792_1;
  assign T_796 = T_794 | T_795;
  assign T_797 = io_tl_acquire_bits_is_builtin_type & T_796;
  assign T_798 = io_tl_acquire_bits_union[11:9];
  assign T_800 = T_797 ? T_798 : 3'h0;
  assign T_801 = {io_tl_acquire_bits_addr_block,io_tl_acquire_bits_addr_beat};
  assign T_802 = {T_801,T_800};
  assign T_803 = io_tl_acquire_bits_union[8:6];
  assign T_813 = 3'h7 == T_803;
  assign T_814 = T_813 ? 3'h3 : 3'h7;
  assign T_815 = 3'h3 == T_803;
  assign T_816 = T_815 ? 3'h3 : T_814;
  assign T_817 = 3'h6 == T_803;
  assign T_818 = T_817 ? 3'h2 : T_816;
  assign T_819 = 3'h2 == T_803;
  assign T_820 = T_819 ? 3'h2 : T_818;
  assign T_821 = 3'h5 == T_803;
  assign T_822 = T_821 ? 3'h1 : T_820;
  assign T_823 = 3'h1 == T_803;
  assign T_824 = T_823 ? 3'h1 : T_822;
  assign T_825 = 3'h4 == T_803;
  assign T_826 = T_825 ? 3'h0 : T_824;
  assign T_827 = 3'h0 == T_803;
  assign T_828 = T_827 ? 3'h0 : T_826;
  assign T_830 = is_subblock ? T_828 : 3'h3;
  assign T_833 = is_subblock ? 3'h0 : 3'h7;
  assign T_853_addr = T_802;
  assign T_853_len = {{5'd0}, T_833};
  assign T_853_size = T_830;
  assign T_853_burst = 2'h1;
  assign T_853_lock = 1'h0;
  assign T_853_cache = 4'h0;
  assign T_853_prot = 3'h0;
  assign T_853_qos = 4'h0;
  assign T_853_region = 4'h0;
  assign T_853_id = get_id_mapper_io_req_out_id;
  assign T_853_user = 1'h0;
  assign T_872 = io_tl_acquire_bits_a_type == 3'h4;
  assign T_873 = io_tl_acquire_bits_is_builtin_type & T_872;
  assign T_875 = T_798[2];
  assign T_877 = 2'h1 << T_875;
  assign T_878 = T_877[0];
  assign T_879 = T_877[1];
  assign T_883 = T_878 ? 4'hf : 4'h0;
  assign T_887 = T_879 ? 4'hf : 4'h0;
  assign T_888 = {T_887,T_883};
  assign T_890 = io_tl_acquire_bits_a_type == 3'h3;
  assign T_891 = io_tl_acquire_bits_is_builtin_type & T_890;
  assign T_893 = io_tl_acquire_bits_a_type == 3'h2;
  assign T_894 = io_tl_acquire_bits_is_builtin_type & T_893;
  assign T_895 = T_891 | T_894;
  assign T_896 = io_tl_acquire_bits_union[8:1];
  assign T_898 = T_895 ? T_896 : 8'h0;
  assign T_899 = T_873 ? T_888 : T_898;
  assign T_900 = ~ T_899;
  assign T_901 = T_900[0];
  assign T_902 = T_900[1];
  assign T_903 = T_900[2];
  assign T_904 = T_900[3];
  assign T_905 = T_900[4];
  assign T_906 = T_900[5];
  assign T_907 = T_900[6];
  assign T_908 = T_900[7];
  assign T_909 = T_901 & T_902;
  assign T_910 = T_903 & T_904;
  assign T_911 = T_905 & T_906;
  assign T_912 = T_907 & T_908;
  assign T_913 = T_909 & T_910;
  assign T_914 = T_911 & T_912;
  assign T_921 = T_914 | T_913;
  assign T_922 = {1'h0,T_913};
  assign T_924 = T_921 ? 2'h2 : 2'h3;
  assign T_925 = T_914 & T_910;
  assign T_926 = T_914 & T_909;
  assign T_927 = T_913 & T_912;
  assign T_928 = T_913 & T_911;
  assign T_929 = T_926 | T_928;
  assign T_930 = T_925 | T_926;
  assign T_931 = T_930 | T_927;
  assign T_932 = T_931 | T_928;
  assign T_933 = {T_922,T_929};
  assign T_935 = T_932 ? 2'h1 : T_924;
  assign T_936 = T_925 & T_902;
  assign T_937 = T_925 & T_901;
  assign T_938 = T_926 & T_904;
  assign T_939 = T_926 & T_903;
  assign T_940 = T_927 & T_906;
  assign T_941 = T_927 & T_905;
  assign T_942 = T_928 & T_908;
  assign T_943 = T_928 & T_907;
  assign T_944 = T_937 | T_939;
  assign T_945 = T_944 | T_941;
  assign T_946 = T_945 | T_943;
  assign T_947 = T_936 | T_937;
  assign T_948 = T_947 | T_938;
  assign T_949 = T_948 | T_939;
  assign T_950 = T_949 | T_940;
  assign T_951 = T_950 | T_941;
  assign T_952 = T_951 | T_942;
  assign T_953 = T_952 | T_943;
  assign put_offset = {T_933,T_946};
  assign put_size = T_953 ? 2'h0 : T_935;
  assign T_956 = w_inflight == 1'h0;
  assign T_957 = put_valid & io_nasti_w_ready;
  assign T_958 = T_957 & put_id_ready;
  assign T_959 = T_958 & T_956;
  assign T_967_0 = 3'h0;
  assign T_967_1 = 3'h4;
  assign T_969 = io_tl_acquire_bits_a_type == T_967_0;
  assign T_970 = io_tl_acquire_bits_a_type == T_967_1;
  assign T_971 = T_969 | T_970;
  assign T_972 = io_tl_acquire_bits_is_builtin_type & T_971;
  assign T_975 = T_972 ? T_798 : 3'h0;
  assign T_977 = {T_801,T_975};
  assign T_979 = is_multibeat ? 4'h0 : put_offset;
  assign GEN_7 = {{28'd0}, T_979};
  assign T_980 = T_977 | GEN_7;
  assign T_982 = is_multibeat ? 2'h3 : put_size;
  assign T_985 = is_multibeat ? 3'h7 : 3'h0;
  assign T_998_addr = T_980;
  assign T_998_len = {{5'd0}, T_985};
  assign T_998_size = {{1'd0}, T_982};
  assign T_998_burst = 2'h1;
  assign T_998_lock = 1'h0;
  assign T_998_cache = 4'h0;
  assign T_998_prot = 3'h0;
  assign T_998_qos = 4'h0;
  assign T_998_region = 4'h0;
  assign T_998_id = put_id_mapper_io_req_out_id;
  assign T_998_user = 1'h0;
  assign T_1017 = T_779 & put_id_ready;
  assign T_1050 = is_multibeat == 1'h0;
  assign T_1051 = w_inflight ? T_725 : T_1050;
  assign T_1058_data = io_tl_acquire_bits_data;
  assign T_1058_last = T_1051;
  assign T_1058_id = w_id;
  assign T_1058_strb = T_899;
  assign T_1058_user = 1'h0;
  assign T_1065 = aw_ready & io_nasti_w_ready;
  assign T_1066 = T_1065 & put_id_ready;
  assign T_1067 = roq_io_enq_ready & io_nasti_ar_ready;
  assign T_1068 = T_1067 & get_id_mapper_io_req_ready;
  assign T_1069 = has_data ? T_1066 : T_1068;
  assign T_1073 = T_956 & T_721;
  assign T_1074 = T_1073 & is_multibeat;
  assign GEN_2 = T_1074 ? 1'h1 : w_inflight;
  assign GEN_3 = T_1074 ? put_id_mapper_io_req_out_id : w_id;
  assign GEN_4 = tl_wrap_out ? 1'h0 : GEN_2;
  assign GEN_5 = w_inflight ? GEN_4 : GEN_2;
  assign T_1077 = io_tl_grant_ready & io_tl_grant_valid;
  assign T_1085_0 = 3'h5;
  assign GEN_8 = {{1'd0}, T_1085_0};
  assign T_1087 = io_tl_grant_bits_g_type == GEN_8;
  assign T_1088 = io_tl_grant_bits_g_type == 4'h0;
  assign T_1089 = io_tl_grant_bits_is_builtin_type ? T_1087 : T_1088;
  assign T_1091 = T_1077 & T_1089;
  assign T_1096 = tl_cnt_in + 3'h1;
  assign T_1097 = T_1096[2:0];
  assign GEN_6 = T_1091 ? T_1097 : tl_cnt_in;
  assign gnt_arb_clk = clk;
  assign gnt_arb_reset = reset;
  assign gnt_arb_io_in_0_valid = io_nasti_r_valid;
  assign gnt_arb_io_in_0_bits_addr_beat = T_1159_addr_beat;
  assign gnt_arb_io_in_0_bits_client_xact_id = T_1159_client_xact_id;
  assign gnt_arb_io_in_0_bits_manager_xact_id = T_1159_manager_xact_id;
  assign gnt_arb_io_in_0_bits_is_builtin_type = T_1159_is_builtin_type;
  assign gnt_arb_io_in_0_bits_g_type = T_1159_g_type;
  assign gnt_arb_io_in_0_bits_data = T_1159_data;
  assign gnt_arb_io_in_0_bits_client_id = GEN_9;
  assign gnt_arb_io_in_1_valid = io_nasti_b_valid;
  assign gnt_arb_io_in_1_bits_addr_beat = T_1230_addr_beat;
  assign gnt_arb_io_in_1_bits_client_xact_id = T_1230_client_xact_id;
  assign gnt_arb_io_in_1_bits_manager_xact_id = T_1230_manager_xact_id;
  assign gnt_arb_io_in_1_bits_is_builtin_type = T_1230_is_builtin_type;
  assign gnt_arb_io_in_1_bits_g_type = T_1230_g_type;
  assign gnt_arb_io_in_1_bits_data = T_1230_data;
  assign gnt_arb_io_in_1_bits_client_id = GEN_10;
  assign gnt_arb_io_out_ready = io_tl_grant_ready;
  assign T_1129 = roq_io_deq_data_subblock ? 3'h4 : 3'h5;
  assign T_1131 = roq_io_deq_data_subblock ? roq_io_deq_data_addr_beat : tl_cnt_in;
  assign T_1159_addr_beat = T_1131;
  assign T_1159_client_xact_id = get_id_mapper_io_resp_in_id;
  assign T_1159_manager_xact_id = 1'h0;
  assign T_1159_is_builtin_type = 1'h1;
  assign T_1159_g_type = {{1'd0}, T_1129};
  assign T_1159_data = io_nasti_r_bits_data;
  assign T_1187 = roq_io_deq_valid == 1'h0;
  assign T_1188 = T_1187 | roq_io_deq_matches;
  assign T_1189 = T_1188 | reset;
  assign T_1191 = T_1189 == 1'h0;
  assign T_1193 = gnt_arb_io_in_0_valid == 1'h0;
  assign T_1194 = T_1193 | get_id_mapper_io_resp_matches;
  assign T_1195 = T_1194 | reset;
  assign T_1197 = T_1195 == 1'h0;
  assign T_1230_addr_beat = 3'h0;
  assign T_1230_client_xact_id = put_id_mapper_io_resp_in_id;
  assign T_1230_manager_xact_id = 1'h0;
  assign T_1230_is_builtin_type = 1'h1;
  assign T_1230_g_type = 4'h3;
  assign T_1230_data = 64'h0;
  assign T_1258 = gnt_arb_io_in_1_valid == 1'h0;
  assign T_1259 = T_1258 | put_id_mapper_io_resp_matches;
  assign T_1260 = T_1259 | reset;
  assign T_1262 = T_1260 == 1'h0;
  assign T_1264 = io_nasti_r_valid == 1'h0;
  assign T_1266 = io_nasti_r_bits_resp == 2'h0;
  assign T_1267 = T_1264 | T_1266;
  assign T_1268 = T_1267 | reset;
  assign T_1270 = T_1268 == 1'h0;
  assign T_1272 = io_nasti_b_valid == 1'h0;
  assign T_1274 = io_nasti_b_bits_resp == 2'h0;
  assign T_1275 = T_1272 | T_1274;
  assign T_1276 = T_1275 | reset;
  assign T_1278 = T_1276 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_11 = {1{$random}};
  tl_cnt_out = GEN_11[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_12 = {1{$random}};
  w_inflight = GEN_12[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_13 = {1{$random}};
  w_id = GEN_13[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_14 = {1{$random}};
  nasti_cnt_out = GEN_14[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_15 = {1{$random}};
  tl_cnt_in = GEN_15[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_16 = {1{$random}};
  GEN_9 = GEN_16[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_17 = {1{$random}};
  GEN_10 = GEN_17[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      tl_cnt_out <= 3'h0;
    end else begin
      if(T_722) begin
        tl_cnt_out <= T_728;
      end
    end
    if(reset) begin
      w_inflight <= 1'h0;
    end else begin
      if(w_inflight) begin
        if(tl_wrap_out) begin
          w_inflight <= 1'h0;
        end else begin
          if(T_1074) begin
            w_inflight <= 1'h1;
          end
        end
      end else begin
        if(T_1074) begin
          w_inflight <= 1'h1;
        end
      end
    end
    if(reset) begin
      w_id <= 5'h0;
    end else begin
      if(T_1074) begin
        w_id <= put_id_mapper_io_req_out_id;
      end
    end
    if(reset) begin
      nasti_cnt_out <= 3'h0;
    end else begin
      if(T_763) begin
        nasti_cnt_out <= T_769;
      end
    end
    if(reset) begin
      tl_cnt_in <= 3'h0;
    end else begin
      if(T_1091) begin
        tl_cnt_in <= T_1097;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1191) begin
          $fwrite(32'h80000002,"Assertion failed: TL -> NASTI converter ReorderQueue: NASTI tag error\n    at Nasti.scala:229 assert(!roq.io.deq.valid || roq.io.deq.matches,\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1191) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1197) begin
          $fwrite(32'h80000002,"Assertion failed: TL -> NASTI ID Mapper: NASTI tag error\n    at Nasti.scala:231 assert(!gnt_arb.io.in(0).valid || get_id_mapper.io.resp.matches,\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1197) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1262) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI tag error\n    at Nasti.scala:243 assert(!gnt_arb.io.in(1).valid || put_id_mapper.io.resp.matches, ---NASTI tag error---)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1262) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1270) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI read error\n    at Nasti.scala:245 assert(!io.nasti.r.valid || io.nasti.r.bits.resp === UInt(0), ---NASTI read error---)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1270) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1278) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI write error\n    at Nasti.scala:246 assert(!io.nasti.b.valid || io.nasti.b.bits.resp === UInt(0), ---NASTI write error---)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1278) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module Queue_10(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [31:0] io_enq_bits_addr,
  input  [7:0] io_enq_bits_len,
  input  [2:0] io_enq_bits_size,
  input  [1:0] io_enq_bits_burst,
  input   io_enq_bits_lock,
  input  [3:0] io_enq_bits_cache,
  input  [2:0] io_enq_bits_prot,
  input  [3:0] io_enq_bits_qos,
  input  [3:0] io_enq_bits_region,
  input  [4:0] io_enq_bits_id,
  input   io_enq_bits_user,
  input   io_deq_ready,
  output  io_deq_valid,
  output [31:0] io_deq_bits_addr,
  output [7:0] io_deq_bits_len,
  output [2:0] io_deq_bits_size,
  output [1:0] io_deq_bits_burst,
  output  io_deq_bits_lock,
  output [3:0] io_deq_bits_cache,
  output [2:0] io_deq_bits_prot,
  output [3:0] io_deq_bits_qos,
  output [3:0] io_deq_bits_region,
  output [4:0] io_deq_bits_id,
  output  io_deq_bits_user,
  output  io_count
);
  reg [31:0] ram_addr [0:0];
  reg [31:0] GEN_0;
  wire [31:0] ram_addr_T_144_data;
  wire  ram_addr_T_144_addr;
  wire  ram_addr_T_144_en;
  wire [31:0] ram_addr_T_125_data;
  wire  ram_addr_T_125_addr;
  wire  ram_addr_T_125_mask;
  wire  ram_addr_T_125_en;
  reg [7:0] ram_len [0:0];
  reg [31:0] GEN_1;
  wire [7:0] ram_len_T_144_data;
  wire  ram_len_T_144_addr;
  wire  ram_len_T_144_en;
  wire [7:0] ram_len_T_125_data;
  wire  ram_len_T_125_addr;
  wire  ram_len_T_125_mask;
  wire  ram_len_T_125_en;
  reg [2:0] ram_size [0:0];
  reg [31:0] GEN_2;
  wire [2:0] ram_size_T_144_data;
  wire  ram_size_T_144_addr;
  wire  ram_size_T_144_en;
  wire [2:0] ram_size_T_125_data;
  wire  ram_size_T_125_addr;
  wire  ram_size_T_125_mask;
  wire  ram_size_T_125_en;
  reg [1:0] ram_burst [0:0];
  reg [31:0] GEN_3;
  wire [1:0] ram_burst_T_144_data;
  wire  ram_burst_T_144_addr;
  wire  ram_burst_T_144_en;
  wire [1:0] ram_burst_T_125_data;
  wire  ram_burst_T_125_addr;
  wire  ram_burst_T_125_mask;
  wire  ram_burst_T_125_en;
  reg  ram_lock [0:0];
  reg [31:0] GEN_4;
  wire  ram_lock_T_144_data;
  wire  ram_lock_T_144_addr;
  wire  ram_lock_T_144_en;
  wire  ram_lock_T_125_data;
  wire  ram_lock_T_125_addr;
  wire  ram_lock_T_125_mask;
  wire  ram_lock_T_125_en;
  reg [3:0] ram_cache [0:0];
  reg [31:0] GEN_5;
  wire [3:0] ram_cache_T_144_data;
  wire  ram_cache_T_144_addr;
  wire  ram_cache_T_144_en;
  wire [3:0] ram_cache_T_125_data;
  wire  ram_cache_T_125_addr;
  wire  ram_cache_T_125_mask;
  wire  ram_cache_T_125_en;
  reg [2:0] ram_prot [0:0];
  reg [31:0] GEN_6;
  wire [2:0] ram_prot_T_144_data;
  wire  ram_prot_T_144_addr;
  wire  ram_prot_T_144_en;
  wire [2:0] ram_prot_T_125_data;
  wire  ram_prot_T_125_addr;
  wire  ram_prot_T_125_mask;
  wire  ram_prot_T_125_en;
  reg [3:0] ram_qos [0:0];
  reg [31:0] GEN_7;
  wire [3:0] ram_qos_T_144_data;
  wire  ram_qos_T_144_addr;
  wire  ram_qos_T_144_en;
  wire [3:0] ram_qos_T_125_data;
  wire  ram_qos_T_125_addr;
  wire  ram_qos_T_125_mask;
  wire  ram_qos_T_125_en;
  reg [3:0] ram_region [0:0];
  reg [31:0] GEN_8;
  wire [3:0] ram_region_T_144_data;
  wire  ram_region_T_144_addr;
  wire  ram_region_T_144_en;
  wire [3:0] ram_region_T_125_data;
  wire  ram_region_T_125_addr;
  wire  ram_region_T_125_mask;
  wire  ram_region_T_125_en;
  reg [4:0] ram_id [0:0];
  reg [31:0] GEN_9;
  wire [4:0] ram_id_T_144_data;
  wire  ram_id_T_144_addr;
  wire  ram_id_T_144_en;
  wire [4:0] ram_id_T_125_data;
  wire  ram_id_T_125_addr;
  wire  ram_id_T_125_mask;
  wire  ram_id_T_125_en;
  reg  ram_user [0:0];
  reg [31:0] GEN_10;
  wire  ram_user_T_144_data;
  wire  ram_user_T_144_addr;
  wire  ram_user_T_144_en;
  wire  ram_user_T_125_data;
  wire  ram_user_T_125_addr;
  wire  ram_user_T_125_mask;
  wire  ram_user_T_125_en;
  reg  maybe_full;
  reg [31:0] GEN_11;
  wire  T_122;
  wire  T_123;
  wire  do_enq;
  wire  T_124;
  wire  do_deq;
  wire  T_139;
  wire  GEN_25;
  wire  T_141;
  wire [1:0] T_156;
  wire  ptr_diff;
  wire [1:0] T_158;
  assign io_enq_ready = T_122;
  assign io_deq_valid = T_141;
  assign io_deq_bits_addr = ram_addr_T_144_data;
  assign io_deq_bits_len = ram_len_T_144_data;
  assign io_deq_bits_size = ram_size_T_144_data;
  assign io_deq_bits_burst = ram_burst_T_144_data;
  assign io_deq_bits_lock = ram_lock_T_144_data;
  assign io_deq_bits_cache = ram_cache_T_144_data;
  assign io_deq_bits_prot = ram_prot_T_144_data;
  assign io_deq_bits_qos = ram_qos_T_144_data;
  assign io_deq_bits_region = ram_region_T_144_data;
  assign io_deq_bits_id = ram_id_T_144_data;
  assign io_deq_bits_user = ram_user_T_144_data;
  assign io_count = T_158[0];
  assign ram_addr_T_144_addr = 1'h0;
  assign ram_addr_T_144_en = 1'h1;
  assign ram_addr_T_144_data = ram_addr[ram_addr_T_144_addr];
  assign ram_addr_T_125_data = io_enq_bits_addr;
  assign ram_addr_T_125_addr = 1'h0;
  assign ram_addr_T_125_mask = do_enq;
  assign ram_addr_T_125_en = do_enq;
  assign ram_len_T_144_addr = 1'h0;
  assign ram_len_T_144_en = 1'h1;
  assign ram_len_T_144_data = ram_len[ram_len_T_144_addr];
  assign ram_len_T_125_data = io_enq_bits_len;
  assign ram_len_T_125_addr = 1'h0;
  assign ram_len_T_125_mask = do_enq;
  assign ram_len_T_125_en = do_enq;
  assign ram_size_T_144_addr = 1'h0;
  assign ram_size_T_144_en = 1'h1;
  assign ram_size_T_144_data = ram_size[ram_size_T_144_addr];
  assign ram_size_T_125_data = io_enq_bits_size;
  assign ram_size_T_125_addr = 1'h0;
  assign ram_size_T_125_mask = do_enq;
  assign ram_size_T_125_en = do_enq;
  assign ram_burst_T_144_addr = 1'h0;
  assign ram_burst_T_144_en = 1'h1;
  assign ram_burst_T_144_data = ram_burst[ram_burst_T_144_addr];
  assign ram_burst_T_125_data = io_enq_bits_burst;
  assign ram_burst_T_125_addr = 1'h0;
  assign ram_burst_T_125_mask = do_enq;
  assign ram_burst_T_125_en = do_enq;
  assign ram_lock_T_144_addr = 1'h0;
  assign ram_lock_T_144_en = 1'h1;
  assign ram_lock_T_144_data = ram_lock[ram_lock_T_144_addr];
  assign ram_lock_T_125_data = io_enq_bits_lock;
  assign ram_lock_T_125_addr = 1'h0;
  assign ram_lock_T_125_mask = do_enq;
  assign ram_lock_T_125_en = do_enq;
  assign ram_cache_T_144_addr = 1'h0;
  assign ram_cache_T_144_en = 1'h1;
  assign ram_cache_T_144_data = ram_cache[ram_cache_T_144_addr];
  assign ram_cache_T_125_data = io_enq_bits_cache;
  assign ram_cache_T_125_addr = 1'h0;
  assign ram_cache_T_125_mask = do_enq;
  assign ram_cache_T_125_en = do_enq;
  assign ram_prot_T_144_addr = 1'h0;
  assign ram_prot_T_144_en = 1'h1;
  assign ram_prot_T_144_data = ram_prot[ram_prot_T_144_addr];
  assign ram_prot_T_125_data = io_enq_bits_prot;
  assign ram_prot_T_125_addr = 1'h0;
  assign ram_prot_T_125_mask = do_enq;
  assign ram_prot_T_125_en = do_enq;
  assign ram_qos_T_144_addr = 1'h0;
  assign ram_qos_T_144_en = 1'h1;
  assign ram_qos_T_144_data = ram_qos[ram_qos_T_144_addr];
  assign ram_qos_T_125_data = io_enq_bits_qos;
  assign ram_qos_T_125_addr = 1'h0;
  assign ram_qos_T_125_mask = do_enq;
  assign ram_qos_T_125_en = do_enq;
  assign ram_region_T_144_addr = 1'h0;
  assign ram_region_T_144_en = 1'h1;
  assign ram_region_T_144_data = ram_region[ram_region_T_144_addr];
  assign ram_region_T_125_data = io_enq_bits_region;
  assign ram_region_T_125_addr = 1'h0;
  assign ram_region_T_125_mask = do_enq;
  assign ram_region_T_125_en = do_enq;
  assign ram_id_T_144_addr = 1'h0;
  assign ram_id_T_144_en = 1'h1;
  assign ram_id_T_144_data = ram_id[ram_id_T_144_addr];
  assign ram_id_T_125_data = io_enq_bits_id;
  assign ram_id_T_125_addr = 1'h0;
  assign ram_id_T_125_mask = do_enq;
  assign ram_id_T_125_en = do_enq;
  assign ram_user_T_144_addr = 1'h0;
  assign ram_user_T_144_en = 1'h1;
  assign ram_user_T_144_data = ram_user[ram_user_T_144_addr];
  assign ram_user_T_125_data = io_enq_bits_user;
  assign ram_user_T_125_addr = 1'h0;
  assign ram_user_T_125_mask = do_enq;
  assign ram_user_T_125_en = do_enq;
  assign T_122 = maybe_full == 1'h0;
  assign T_123 = io_enq_ready & io_enq_valid;
  assign do_enq = T_123;
  assign T_124 = io_deq_ready & io_deq_valid;
  assign do_deq = T_124;
  assign T_139 = do_enq != do_deq;
  assign GEN_25 = T_139 ? do_enq : maybe_full;
  assign T_141 = T_122 == 1'h0;
  assign T_156 = 1'h0 - 1'h0;
  assign ptr_diff = T_156[0:0];
  assign T_158 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = GEN_0[31:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = GEN_1[7:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = GEN_2[2:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_burst[initvar] = GEN_3[1:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_lock[initvar] = GEN_4[0:0];
  `endif
  GEN_5 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_cache[initvar] = GEN_5[3:0];
  `endif
  GEN_6 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_prot[initvar] = GEN_6[2:0];
  `endif
  GEN_7 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_qos[initvar] = GEN_7[3:0];
  `endif
  GEN_8 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_region[initvar] = GEN_8[3:0];
  `endif
  GEN_9 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = GEN_9[4:0];
  `endif
  GEN_10 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_user[initvar] = GEN_10[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_11 = {1{$random}};
  maybe_full = GEN_11[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_addr_T_125_en & ram_addr_T_125_mask) begin
      ram_addr[ram_addr_T_125_addr] <= ram_addr_T_125_data;
    end
    if(ram_len_T_125_en & ram_len_T_125_mask) begin
      ram_len[ram_len_T_125_addr] <= ram_len_T_125_data;
    end
    if(ram_size_T_125_en & ram_size_T_125_mask) begin
      ram_size[ram_size_T_125_addr] <= ram_size_T_125_data;
    end
    if(ram_burst_T_125_en & ram_burst_T_125_mask) begin
      ram_burst[ram_burst_T_125_addr] <= ram_burst_T_125_data;
    end
    if(ram_lock_T_125_en & ram_lock_T_125_mask) begin
      ram_lock[ram_lock_T_125_addr] <= ram_lock_T_125_data;
    end
    if(ram_cache_T_125_en & ram_cache_T_125_mask) begin
      ram_cache[ram_cache_T_125_addr] <= ram_cache_T_125_data;
    end
    if(ram_prot_T_125_en & ram_prot_T_125_mask) begin
      ram_prot[ram_prot_T_125_addr] <= ram_prot_T_125_data;
    end
    if(ram_qos_T_125_en & ram_qos_T_125_mask) begin
      ram_qos[ram_qos_T_125_addr] <= ram_qos_T_125_data;
    end
    if(ram_region_T_125_en & ram_region_T_125_mask) begin
      ram_region[ram_region_T_125_addr] <= ram_region_T_125_data;
    end
    if(ram_id_T_125_en & ram_id_T_125_mask) begin
      ram_id[ram_id_T_125_addr] <= ram_id_T_125_data;
    end
    if(ram_user_T_125_en & ram_user_T_125_mask) begin
      ram_user[ram_user_T_125_addr] <= ram_user_T_125_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_139) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_12(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [63:0] io_enq_bits_data,
  input   io_enq_bits_last,
  input  [4:0] io_enq_bits_id,
  input  [7:0] io_enq_bits_strb,
  input   io_enq_bits_user,
  input   io_deq_ready,
  output  io_deq_valid,
  output [63:0] io_deq_bits_data,
  output  io_deq_bits_last,
  output [4:0] io_deq_bits_id,
  output [7:0] io_deq_bits_strb,
  output  io_deq_bits_user,
  output [1:0] io_count
);
  reg [63:0] ram_data [0:1];
  reg [63:0] GEN_0;
  wire [63:0] ram_data_T_94_data;
  wire  ram_data_T_94_addr;
  wire  ram_data_T_94_en;
  wire [63:0] ram_data_T_73_data;
  wire  ram_data_T_73_addr;
  wire  ram_data_T_73_mask;
  wire  ram_data_T_73_en;
  reg  ram_last [0:1];
  reg [31:0] GEN_1;
  wire  ram_last_T_94_data;
  wire  ram_last_T_94_addr;
  wire  ram_last_T_94_en;
  wire  ram_last_T_73_data;
  wire  ram_last_T_73_addr;
  wire  ram_last_T_73_mask;
  wire  ram_last_T_73_en;
  reg [4:0] ram_id [0:1];
  reg [31:0] GEN_2;
  wire [4:0] ram_id_T_94_data;
  wire  ram_id_T_94_addr;
  wire  ram_id_T_94_en;
  wire [4:0] ram_id_T_73_data;
  wire  ram_id_T_73_addr;
  wire  ram_id_T_73_mask;
  wire  ram_id_T_73_en;
  reg [7:0] ram_strb [0:1];
  reg [31:0] GEN_3;
  wire [7:0] ram_strb_T_94_data;
  wire  ram_strb_T_94_addr;
  wire  ram_strb_T_94_en;
  wire [7:0] ram_strb_T_73_data;
  wire  ram_strb_T_73_addr;
  wire  ram_strb_T_73_mask;
  wire  ram_strb_T_73_en;
  reg  ram_user [0:1];
  reg [31:0] GEN_4;
  wire  ram_user_T_94_data;
  wire  ram_user_T_94_addr;
  wire  ram_user_T_94_en;
  wire  ram_user_T_73_data;
  wire  ram_user_T_73_addr;
  wire  ram_user_T_73_mask;
  wire  ram_user_T_73_en;
  reg  T_65;
  reg [31:0] GEN_5;
  reg  T_67;
  reg [31:0] GEN_6;
  reg  maybe_full;
  reg [31:0] GEN_7;
  wire  ptr_match;
  wire  T_70;
  wire  empty;
  wire  full;
  wire  T_71;
  wire  do_enq;
  wire  T_72;
  wire  do_deq;
  wire [1:0] T_82;
  wire  T_83;
  wire  GEN_13;
  wire [1:0] T_87;
  wire  T_88;
  wire  GEN_14;
  wire  T_89;
  wire  GEN_15;
  wire  T_91;
  wire  T_93;
  wire [1:0] T_100;
  wire  ptr_diff;
  wire  T_101;
  wire [1:0] T_102;
  assign io_enq_ready = T_93;
  assign io_deq_valid = T_91;
  assign io_deq_bits_data = ram_data_T_94_data;
  assign io_deq_bits_last = ram_last_T_94_data;
  assign io_deq_bits_id = ram_id_T_94_data;
  assign io_deq_bits_strb = ram_strb_T_94_data;
  assign io_deq_bits_user = ram_user_T_94_data;
  assign io_count = T_102;
  assign ram_data_T_94_addr = T_67;
  assign ram_data_T_94_en = 1'h1;
  assign ram_data_T_94_data = ram_data[ram_data_T_94_addr];
  assign ram_data_T_73_data = io_enq_bits_data;
  assign ram_data_T_73_addr = T_65;
  assign ram_data_T_73_mask = do_enq;
  assign ram_data_T_73_en = do_enq;
  assign ram_last_T_94_addr = T_67;
  assign ram_last_T_94_en = 1'h1;
  assign ram_last_T_94_data = ram_last[ram_last_T_94_addr];
  assign ram_last_T_73_data = io_enq_bits_last;
  assign ram_last_T_73_addr = T_65;
  assign ram_last_T_73_mask = do_enq;
  assign ram_last_T_73_en = do_enq;
  assign ram_id_T_94_addr = T_67;
  assign ram_id_T_94_en = 1'h1;
  assign ram_id_T_94_data = ram_id[ram_id_T_94_addr];
  assign ram_id_T_73_data = io_enq_bits_id;
  assign ram_id_T_73_addr = T_65;
  assign ram_id_T_73_mask = do_enq;
  assign ram_id_T_73_en = do_enq;
  assign ram_strb_T_94_addr = T_67;
  assign ram_strb_T_94_en = 1'h1;
  assign ram_strb_T_94_data = ram_strb[ram_strb_T_94_addr];
  assign ram_strb_T_73_data = io_enq_bits_strb;
  assign ram_strb_T_73_addr = T_65;
  assign ram_strb_T_73_mask = do_enq;
  assign ram_strb_T_73_en = do_enq;
  assign ram_user_T_94_addr = T_67;
  assign ram_user_T_94_en = 1'h1;
  assign ram_user_T_94_data = ram_user[ram_user_T_94_addr];
  assign ram_user_T_73_data = io_enq_bits_user;
  assign ram_user_T_73_addr = T_65;
  assign ram_user_T_73_mask = do_enq;
  assign ram_user_T_73_en = do_enq;
  assign ptr_match = T_65 == T_67;
  assign T_70 = maybe_full == 1'h0;
  assign empty = ptr_match & T_70;
  assign full = ptr_match & maybe_full;
  assign T_71 = io_enq_ready & io_enq_valid;
  assign do_enq = T_71;
  assign T_72 = io_deq_ready & io_deq_valid;
  assign do_deq = T_72;
  assign T_82 = T_65 + 1'h1;
  assign T_83 = T_82[0:0];
  assign GEN_13 = do_enq ? T_83 : T_65;
  assign T_87 = T_67 + 1'h1;
  assign T_88 = T_87[0:0];
  assign GEN_14 = do_deq ? T_88 : T_67;
  assign T_89 = do_enq != do_deq;
  assign GEN_15 = T_89 ? do_enq : maybe_full;
  assign T_91 = empty == 1'h0;
  assign T_93 = full == 1'h0;
  assign T_100 = T_65 - T_67;
  assign ptr_diff = T_100[0:0];
  assign T_101 = maybe_full & ptr_match;
  assign T_102 = {T_101,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {2{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = GEN_0[63:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_last[initvar] = GEN_1[0:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = GEN_2[4:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_strb[initvar] = GEN_3[7:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user[initvar] = GEN_4[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_5 = {1{$random}};
  T_65 = GEN_5[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_6 = {1{$random}};
  T_67 = GEN_6[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_7 = {1{$random}};
  maybe_full = GEN_7[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_data_T_73_en & ram_data_T_73_mask) begin
      ram_data[ram_data_T_73_addr] <= ram_data_T_73_data;
    end
    if(ram_last_T_73_en & ram_last_T_73_mask) begin
      ram_last[ram_last_T_73_addr] <= ram_last_T_73_data;
    end
    if(ram_id_T_73_en & ram_id_T_73_mask) begin
      ram_id[ram_id_T_73_addr] <= ram_id_T_73_data;
    end
    if(ram_strb_T_73_en & ram_strb_T_73_mask) begin
      ram_strb[ram_strb_T_73_addr] <= ram_strb_T_73_data;
    end
    if(ram_user_T_73_en & ram_user_T_73_mask) begin
      ram_user[ram_user_T_73_addr] <= ram_user_T_73_data;
    end
    if(reset) begin
      T_65 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_65 <= T_83;
      end
    end
    if(reset) begin
      T_67 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_67 <= T_88;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_89) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_13(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_resp,
  input  [63:0] io_enq_bits_data,
  input   io_enq_bits_last,
  input  [4:0] io_enq_bits_id,
  input   io_enq_bits_user,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_resp,
  output [63:0] io_deq_bits_data,
  output  io_deq_bits_last,
  output [4:0] io_deq_bits_id,
  output  io_deq_bits_user,
  output [1:0] io_count
);
  reg [1:0] ram_resp [0:1];
  reg [31:0] GEN_0;
  wire [1:0] ram_resp_T_94_data;
  wire  ram_resp_T_94_addr;
  wire  ram_resp_T_94_en;
  wire [1:0] ram_resp_T_73_data;
  wire  ram_resp_T_73_addr;
  wire  ram_resp_T_73_mask;
  wire  ram_resp_T_73_en;
  reg [63:0] ram_data [0:1];
  reg [63:0] GEN_1;
  wire [63:0] ram_data_T_94_data;
  wire  ram_data_T_94_addr;
  wire  ram_data_T_94_en;
  wire [63:0] ram_data_T_73_data;
  wire  ram_data_T_73_addr;
  wire  ram_data_T_73_mask;
  wire  ram_data_T_73_en;
  reg  ram_last [0:1];
  reg [31:0] GEN_2;
  wire  ram_last_T_94_data;
  wire  ram_last_T_94_addr;
  wire  ram_last_T_94_en;
  wire  ram_last_T_73_data;
  wire  ram_last_T_73_addr;
  wire  ram_last_T_73_mask;
  wire  ram_last_T_73_en;
  reg [4:0] ram_id [0:1];
  reg [31:0] GEN_3;
  wire [4:0] ram_id_T_94_data;
  wire  ram_id_T_94_addr;
  wire  ram_id_T_94_en;
  wire [4:0] ram_id_T_73_data;
  wire  ram_id_T_73_addr;
  wire  ram_id_T_73_mask;
  wire  ram_id_T_73_en;
  reg  ram_user [0:1];
  reg [31:0] GEN_4;
  wire  ram_user_T_94_data;
  wire  ram_user_T_94_addr;
  wire  ram_user_T_94_en;
  wire  ram_user_T_73_data;
  wire  ram_user_T_73_addr;
  wire  ram_user_T_73_mask;
  wire  ram_user_T_73_en;
  reg  T_65;
  reg [31:0] GEN_5;
  reg  T_67;
  reg [31:0] GEN_6;
  reg  maybe_full;
  reg [31:0] GEN_7;
  wire  ptr_match;
  wire  T_70;
  wire  empty;
  wire  full;
  wire  T_71;
  wire  do_enq;
  wire  T_72;
  wire  do_deq;
  wire [1:0] T_82;
  wire  T_83;
  wire  GEN_13;
  wire [1:0] T_87;
  wire  T_88;
  wire  GEN_14;
  wire  T_89;
  wire  GEN_15;
  wire  T_91;
  wire  T_93;
  wire [1:0] T_100;
  wire  ptr_diff;
  wire  T_101;
  wire [1:0] T_102;
  assign io_enq_ready = T_93;
  assign io_deq_valid = T_91;
  assign io_deq_bits_resp = ram_resp_T_94_data;
  assign io_deq_bits_data = ram_data_T_94_data;
  assign io_deq_bits_last = ram_last_T_94_data;
  assign io_deq_bits_id = ram_id_T_94_data;
  assign io_deq_bits_user = ram_user_T_94_data;
  assign io_count = T_102;
  assign ram_resp_T_94_addr = T_67;
  assign ram_resp_T_94_en = 1'h1;
  assign ram_resp_T_94_data = ram_resp[ram_resp_T_94_addr];
  assign ram_resp_T_73_data = io_enq_bits_resp;
  assign ram_resp_T_73_addr = T_65;
  assign ram_resp_T_73_mask = do_enq;
  assign ram_resp_T_73_en = do_enq;
  assign ram_data_T_94_addr = T_67;
  assign ram_data_T_94_en = 1'h1;
  assign ram_data_T_94_data = ram_data[ram_data_T_94_addr];
  assign ram_data_T_73_data = io_enq_bits_data;
  assign ram_data_T_73_addr = T_65;
  assign ram_data_T_73_mask = do_enq;
  assign ram_data_T_73_en = do_enq;
  assign ram_last_T_94_addr = T_67;
  assign ram_last_T_94_en = 1'h1;
  assign ram_last_T_94_data = ram_last[ram_last_T_94_addr];
  assign ram_last_T_73_data = io_enq_bits_last;
  assign ram_last_T_73_addr = T_65;
  assign ram_last_T_73_mask = do_enq;
  assign ram_last_T_73_en = do_enq;
  assign ram_id_T_94_addr = T_67;
  assign ram_id_T_94_en = 1'h1;
  assign ram_id_T_94_data = ram_id[ram_id_T_94_addr];
  assign ram_id_T_73_data = io_enq_bits_id;
  assign ram_id_T_73_addr = T_65;
  assign ram_id_T_73_mask = do_enq;
  assign ram_id_T_73_en = do_enq;
  assign ram_user_T_94_addr = T_67;
  assign ram_user_T_94_en = 1'h1;
  assign ram_user_T_94_data = ram_user[ram_user_T_94_addr];
  assign ram_user_T_73_data = io_enq_bits_user;
  assign ram_user_T_73_addr = T_65;
  assign ram_user_T_73_mask = do_enq;
  assign ram_user_T_73_en = do_enq;
  assign ptr_match = T_65 == T_67;
  assign T_70 = maybe_full == 1'h0;
  assign empty = ptr_match & T_70;
  assign full = ptr_match & maybe_full;
  assign T_71 = io_enq_ready & io_enq_valid;
  assign do_enq = T_71;
  assign T_72 = io_deq_ready & io_deq_valid;
  assign do_deq = T_72;
  assign T_82 = T_65 + 1'h1;
  assign T_83 = T_82[0:0];
  assign GEN_13 = do_enq ? T_83 : T_65;
  assign T_87 = T_67 + 1'h1;
  assign T_88 = T_87[0:0];
  assign GEN_14 = do_deq ? T_88 : T_67;
  assign T_89 = do_enq != do_deq;
  assign GEN_15 = T_89 ? do_enq : maybe_full;
  assign T_91 = empty == 1'h0;
  assign T_93 = full == 1'h0;
  assign T_100 = T_65 - T_67;
  assign ptr_diff = T_100[0:0];
  assign T_101 = maybe_full & ptr_match;
  assign T_102 = {T_101,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_resp[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {2{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = GEN_1[63:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_last[initvar] = GEN_2[0:0];
  `endif
  GEN_3 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = GEN_3[4:0];
  `endif
  GEN_4 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user[initvar] = GEN_4[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_5 = {1{$random}};
  T_65 = GEN_5[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_6 = {1{$random}};
  T_67 = GEN_6[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_7 = {1{$random}};
  maybe_full = GEN_7[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_resp_T_73_en & ram_resp_T_73_mask) begin
      ram_resp[ram_resp_T_73_addr] <= ram_resp_T_73_data;
    end
    if(ram_data_T_73_en & ram_data_T_73_mask) begin
      ram_data[ram_data_T_73_addr] <= ram_data_T_73_data;
    end
    if(ram_last_T_73_en & ram_last_T_73_mask) begin
      ram_last[ram_last_T_73_addr] <= ram_last_T_73_data;
    end
    if(ram_id_T_73_en & ram_id_T_73_mask) begin
      ram_id[ram_id_T_73_addr] <= ram_id_T_73_data;
    end
    if(ram_user_T_73_en & ram_user_T_73_mask) begin
      ram_user[ram_user_T_73_addr] <= ram_user_T_73_data;
    end
    if(reset) begin
      T_65 <= 1'h0;
    end else begin
      if(do_enq) begin
        T_65 <= T_83;
      end
    end
    if(reset) begin
      T_67 <= 1'h0;
    end else begin
      if(do_deq) begin
        T_67 <= T_88;
      end
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_89) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module Queue_14(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_resp,
  input  [4:0] io_enq_bits_id,
  input   io_enq_bits_user,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_resp,
  output [4:0] io_deq_bits_id,
  output  io_deq_bits_user,
  output  io_count
);
  reg [1:0] ram_resp [0:0];
  reg [31:0] GEN_0;
  wire [1:0] ram_resp_T_64_data;
  wire  ram_resp_T_64_addr;
  wire  ram_resp_T_64_en;
  wire [1:0] ram_resp_T_53_data;
  wire  ram_resp_T_53_addr;
  wire  ram_resp_T_53_mask;
  wire  ram_resp_T_53_en;
  reg [4:0] ram_id [0:0];
  reg [31:0] GEN_1;
  wire [4:0] ram_id_T_64_data;
  wire  ram_id_T_64_addr;
  wire  ram_id_T_64_en;
  wire [4:0] ram_id_T_53_data;
  wire  ram_id_T_53_addr;
  wire  ram_id_T_53_mask;
  wire  ram_id_T_53_en;
  reg  ram_user [0:0];
  reg [31:0] GEN_2;
  wire  ram_user_T_64_data;
  wire  ram_user_T_64_addr;
  wire  ram_user_T_64_en;
  wire  ram_user_T_53_data;
  wire  ram_user_T_53_addr;
  wire  ram_user_T_53_mask;
  wire  ram_user_T_53_en;
  reg  maybe_full;
  reg [31:0] GEN_3;
  wire  T_50;
  wire  T_51;
  wire  do_enq;
  wire  T_52;
  wire  do_deq;
  wire  T_59;
  wire  GEN_9;
  wire  T_61;
  wire [1:0] T_68;
  wire  ptr_diff;
  wire [1:0] T_70;
  assign io_enq_ready = T_50;
  assign io_deq_valid = T_61;
  assign io_deq_bits_resp = ram_resp_T_64_data;
  assign io_deq_bits_id = ram_id_T_64_data;
  assign io_deq_bits_user = ram_user_T_64_data;
  assign io_count = T_70[0];
  assign ram_resp_T_64_addr = 1'h0;
  assign ram_resp_T_64_en = 1'h1;
  assign ram_resp_T_64_data = ram_resp[ram_resp_T_64_addr];
  assign ram_resp_T_53_data = io_enq_bits_resp;
  assign ram_resp_T_53_addr = 1'h0;
  assign ram_resp_T_53_mask = do_enq;
  assign ram_resp_T_53_en = do_enq;
  assign ram_id_T_64_addr = 1'h0;
  assign ram_id_T_64_en = 1'h1;
  assign ram_id_T_64_data = ram_id[ram_id_T_64_addr];
  assign ram_id_T_53_data = io_enq_bits_id;
  assign ram_id_T_53_addr = 1'h0;
  assign ram_id_T_53_mask = do_enq;
  assign ram_id_T_53_en = do_enq;
  assign ram_user_T_64_addr = 1'h0;
  assign ram_user_T_64_en = 1'h1;
  assign ram_user_T_64_data = ram_user[ram_user_T_64_addr];
  assign ram_user_T_53_data = io_enq_bits_user;
  assign ram_user_T_53_addr = 1'h0;
  assign ram_user_T_53_mask = do_enq;
  assign ram_user_T_53_en = do_enq;
  assign T_50 = maybe_full == 1'h0;
  assign T_51 = io_enq_ready & io_enq_valid;
  assign do_enq = T_51;
  assign T_52 = io_deq_ready & io_deq_valid;
  assign do_deq = T_52;
  assign T_59 = do_enq != do_deq;
  assign GEN_9 = T_59 ? do_enq : maybe_full;
  assign T_61 = T_50 == 1'h0;
  assign T_68 = 1'h0 - 1'h0;
  assign ptr_diff = T_68[0:0];
  assign T_70 = {maybe_full,ptr_diff};
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_resp[initvar] = GEN_0[1:0];
  `endif
  GEN_1 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = GEN_1[4:0];
  `endif
  GEN_2 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_user[initvar] = GEN_2[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_3 = {1{$random}};
  maybe_full = GEN_3[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(ram_resp_T_53_en & ram_resp_T_53_mask) begin
      ram_resp[ram_resp_T_53_addr] <= ram_resp_T_53_data;
    end
    if(ram_id_T_53_en & ram_id_T_53_mask) begin
      ram_id[ram_id_T_53_addr] <= ram_id_T_53_data;
    end
    if(ram_user_T_53_en & ram_user_T_53_mask) begin
      ram_user[ram_user_T_53_addr] <= ram_user_T_53_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      if(T_59) begin
        maybe_full <= do_enq;
      end
    end
  end
endmodule
module OuterMemorySystem(
  input   clk,
  input   reset,
  output  io_tiles_cached_0_acquire_ready,
  input   io_tiles_cached_0_acquire_valid,
  input  [25:0] io_tiles_cached_0_acquire_bits_addr_block,
  input   io_tiles_cached_0_acquire_bits_client_xact_id,
  input  [2:0] io_tiles_cached_0_acquire_bits_addr_beat,
  input   io_tiles_cached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_tiles_cached_0_acquire_bits_a_type,
  input  [11:0] io_tiles_cached_0_acquire_bits_union,
  input  [63:0] io_tiles_cached_0_acquire_bits_data,
  input   io_tiles_cached_0_probe_ready,
  output  io_tiles_cached_0_probe_valid,
  output [25:0] io_tiles_cached_0_probe_bits_addr_block,
  output [1:0] io_tiles_cached_0_probe_bits_p_type,
  output  io_tiles_cached_0_release_ready,
  input   io_tiles_cached_0_release_valid,
  input  [2:0] io_tiles_cached_0_release_bits_addr_beat,
  input  [25:0] io_tiles_cached_0_release_bits_addr_block,
  input   io_tiles_cached_0_release_bits_client_xact_id,
  input   io_tiles_cached_0_release_bits_voluntary,
  input  [2:0] io_tiles_cached_0_release_bits_r_type,
  input  [63:0] io_tiles_cached_0_release_bits_data,
  input   io_tiles_cached_0_grant_ready,
  output  io_tiles_cached_0_grant_valid,
  output [2:0] io_tiles_cached_0_grant_bits_addr_beat,
  output  io_tiles_cached_0_grant_bits_client_xact_id,
  output [1:0] io_tiles_cached_0_grant_bits_manager_xact_id,
  output  io_tiles_cached_0_grant_bits_is_builtin_type,
  output [3:0] io_tiles_cached_0_grant_bits_g_type,
  output [63:0] io_tiles_cached_0_grant_bits_data,
  output  io_tiles_cached_0_grant_bits_manager_id,
  output  io_tiles_cached_0_finish_ready,
  input   io_tiles_cached_0_finish_valid,
  input  [1:0] io_tiles_cached_0_finish_bits_manager_xact_id,
  input   io_tiles_cached_0_finish_bits_manager_id,
  output  io_tiles_uncached_0_acquire_ready,
  input   io_tiles_uncached_0_acquire_valid,
  input  [25:0] io_tiles_uncached_0_acquire_bits_addr_block,
  input   io_tiles_uncached_0_acquire_bits_client_xact_id,
  input  [2:0] io_tiles_uncached_0_acquire_bits_addr_beat,
  input   io_tiles_uncached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_tiles_uncached_0_acquire_bits_a_type,
  input  [11:0] io_tiles_uncached_0_acquire_bits_union,
  input  [63:0] io_tiles_uncached_0_acquire_bits_data,
  input   io_tiles_uncached_0_grant_ready,
  output  io_tiles_uncached_0_grant_valid,
  output [2:0] io_tiles_uncached_0_grant_bits_addr_beat,
  output  io_tiles_uncached_0_grant_bits_client_xact_id,
  output [1:0] io_tiles_uncached_0_grant_bits_manager_xact_id,
  output  io_tiles_uncached_0_grant_bits_is_builtin_type,
  output [3:0] io_tiles_uncached_0_grant_bits_g_type,
  output [63:0] io_tiles_uncached_0_grant_bits_data,
  input   io_incoherent_0,
  input   io_mem_axi_0_aw_ready,
  output  io_mem_axi_0_aw_valid,
  output [31:0] io_mem_axi_0_aw_bits_addr,
  output [7:0] io_mem_axi_0_aw_bits_len,
  output [2:0] io_mem_axi_0_aw_bits_size,
  output [1:0] io_mem_axi_0_aw_bits_burst,
  output  io_mem_axi_0_aw_bits_lock,
  output [3:0] io_mem_axi_0_aw_bits_cache,
  output [2:0] io_mem_axi_0_aw_bits_prot,
  output [3:0] io_mem_axi_0_aw_bits_qos,
  output [3:0] io_mem_axi_0_aw_bits_region,
  output [4:0] io_mem_axi_0_aw_bits_id,
  output  io_mem_axi_0_aw_bits_user,
  input   io_mem_axi_0_w_ready,
  output  io_mem_axi_0_w_valid,
  output [63:0] io_mem_axi_0_w_bits_data,
  output  io_mem_axi_0_w_bits_last,
  output [4:0] io_mem_axi_0_w_bits_id,
  output [7:0] io_mem_axi_0_w_bits_strb,
  output  io_mem_axi_0_w_bits_user,
  output  io_mem_axi_0_b_ready,
  input   io_mem_axi_0_b_valid,
  input  [1:0] io_mem_axi_0_b_bits_resp,
  input  [4:0] io_mem_axi_0_b_bits_id,
  input   io_mem_axi_0_b_bits_user,
  input   io_mem_axi_0_ar_ready,
  output  io_mem_axi_0_ar_valid,
  output [31:0] io_mem_axi_0_ar_bits_addr,
  output [7:0] io_mem_axi_0_ar_bits_len,
  output [2:0] io_mem_axi_0_ar_bits_size,
  output [1:0] io_mem_axi_0_ar_bits_burst,
  output  io_mem_axi_0_ar_bits_lock,
  output [3:0] io_mem_axi_0_ar_bits_cache,
  output [2:0] io_mem_axi_0_ar_bits_prot,
  output [3:0] io_mem_axi_0_ar_bits_qos,
  output [3:0] io_mem_axi_0_ar_bits_region,
  output [4:0] io_mem_axi_0_ar_bits_id,
  output  io_mem_axi_0_ar_bits_user,
  output  io_mem_axi_0_r_ready,
  input   io_mem_axi_0_r_valid,
  input  [1:0] io_mem_axi_0_r_bits_resp,
  input  [63:0] io_mem_axi_0_r_bits_data,
  input   io_mem_axi_0_r_bits_last,
  input  [4:0] io_mem_axi_0_r_bits_id,
  input   io_mem_axi_0_r_bits_user,
  input   io_mmio_acquire_ready,
  output  io_mmio_acquire_valid,
  output [25:0] io_mmio_acquire_bits_addr_block,
  output [1:0] io_mmio_acquire_bits_client_xact_id,
  output [2:0] io_mmio_acquire_bits_addr_beat,
  output  io_mmio_acquire_bits_is_builtin_type,
  output [2:0] io_mmio_acquire_bits_a_type,
  output [11:0] io_mmio_acquire_bits_union,
  output [63:0] io_mmio_acquire_bits_data,
  output  io_mmio_grant_ready,
  input   io_mmio_grant_valid,
  input  [2:0] io_mmio_grant_bits_addr_beat,
  input  [1:0] io_mmio_grant_bits_client_xact_id,
  input   io_mmio_grant_bits_manager_xact_id,
  input   io_mmio_grant_bits_is_builtin_type,
  input  [3:0] io_mmio_grant_bits_g_type,
  input  [63:0] io_mmio_grant_bits_data
);
  wire  l1tol2net_clk;
  wire  l1tol2net_reset;
  wire  l1tol2net_io_clients_cached_0_acquire_ready;
  wire  l1tol2net_io_clients_cached_0_acquire_valid;
  wire [25:0] l1tol2net_io_clients_cached_0_acquire_bits_addr_block;
  wire  l1tol2net_io_clients_cached_0_acquire_bits_client_xact_id;
  wire [2:0] l1tol2net_io_clients_cached_0_acquire_bits_addr_beat;
  wire  l1tol2net_io_clients_cached_0_acquire_bits_is_builtin_type;
  wire [2:0] l1tol2net_io_clients_cached_0_acquire_bits_a_type;
  wire [11:0] l1tol2net_io_clients_cached_0_acquire_bits_union;
  wire [63:0] l1tol2net_io_clients_cached_0_acquire_bits_data;
  wire  l1tol2net_io_clients_cached_0_probe_ready;
  wire  l1tol2net_io_clients_cached_0_probe_valid;
  wire [25:0] l1tol2net_io_clients_cached_0_probe_bits_addr_block;
  wire [1:0] l1tol2net_io_clients_cached_0_probe_bits_p_type;
  wire  l1tol2net_io_clients_cached_0_release_ready;
  wire  l1tol2net_io_clients_cached_0_release_valid;
  wire [2:0] l1tol2net_io_clients_cached_0_release_bits_addr_beat;
  wire [25:0] l1tol2net_io_clients_cached_0_release_bits_addr_block;
  wire  l1tol2net_io_clients_cached_0_release_bits_client_xact_id;
  wire  l1tol2net_io_clients_cached_0_release_bits_voluntary;
  wire [2:0] l1tol2net_io_clients_cached_0_release_bits_r_type;
  wire [63:0] l1tol2net_io_clients_cached_0_release_bits_data;
  wire  l1tol2net_io_clients_cached_0_grant_ready;
  wire  l1tol2net_io_clients_cached_0_grant_valid;
  wire [2:0] l1tol2net_io_clients_cached_0_grant_bits_addr_beat;
  wire  l1tol2net_io_clients_cached_0_grant_bits_client_xact_id;
  wire [1:0] l1tol2net_io_clients_cached_0_grant_bits_manager_xact_id;
  wire  l1tol2net_io_clients_cached_0_grant_bits_is_builtin_type;
  wire [3:0] l1tol2net_io_clients_cached_0_grant_bits_g_type;
  wire [63:0] l1tol2net_io_clients_cached_0_grant_bits_data;
  wire  l1tol2net_io_clients_cached_0_grant_bits_manager_id;
  wire  l1tol2net_io_clients_cached_0_finish_ready;
  wire  l1tol2net_io_clients_cached_0_finish_valid;
  wire [1:0] l1tol2net_io_clients_cached_0_finish_bits_manager_xact_id;
  wire  l1tol2net_io_clients_cached_0_finish_bits_manager_id;
  wire  l1tol2net_io_clients_uncached_0_acquire_ready;
  wire  l1tol2net_io_clients_uncached_0_acquire_valid;
  wire [25:0] l1tol2net_io_clients_uncached_0_acquire_bits_addr_block;
  wire  l1tol2net_io_clients_uncached_0_acquire_bits_client_xact_id;
  wire [2:0] l1tol2net_io_clients_uncached_0_acquire_bits_addr_beat;
  wire  l1tol2net_io_clients_uncached_0_acquire_bits_is_builtin_type;
  wire [2:0] l1tol2net_io_clients_uncached_0_acquire_bits_a_type;
  wire [11:0] l1tol2net_io_clients_uncached_0_acquire_bits_union;
  wire [63:0] l1tol2net_io_clients_uncached_0_acquire_bits_data;
  wire  l1tol2net_io_clients_uncached_0_grant_ready;
  wire  l1tol2net_io_clients_uncached_0_grant_valid;
  wire [2:0] l1tol2net_io_clients_uncached_0_grant_bits_addr_beat;
  wire  l1tol2net_io_clients_uncached_0_grant_bits_client_xact_id;
  wire [1:0] l1tol2net_io_clients_uncached_0_grant_bits_manager_xact_id;
  wire  l1tol2net_io_clients_uncached_0_grant_bits_is_builtin_type;
  wire [3:0] l1tol2net_io_clients_uncached_0_grant_bits_g_type;
  wire [63:0] l1tol2net_io_clients_uncached_0_grant_bits_data;
  wire  l1tol2net_io_managers_0_acquire_ready;
  wire  l1tol2net_io_managers_0_acquire_valid;
  wire [25:0] l1tol2net_io_managers_0_acquire_bits_addr_block;
  wire  l1tol2net_io_managers_0_acquire_bits_client_xact_id;
  wire [2:0] l1tol2net_io_managers_0_acquire_bits_addr_beat;
  wire  l1tol2net_io_managers_0_acquire_bits_is_builtin_type;
  wire [2:0] l1tol2net_io_managers_0_acquire_bits_a_type;
  wire [11:0] l1tol2net_io_managers_0_acquire_bits_union;
  wire [63:0] l1tol2net_io_managers_0_acquire_bits_data;
  wire  l1tol2net_io_managers_0_acquire_bits_client_id;
  wire  l1tol2net_io_managers_0_grant_ready;
  wire  l1tol2net_io_managers_0_grant_valid;
  wire [2:0] l1tol2net_io_managers_0_grant_bits_addr_beat;
  wire  l1tol2net_io_managers_0_grant_bits_client_xact_id;
  wire [1:0] l1tol2net_io_managers_0_grant_bits_manager_xact_id;
  wire  l1tol2net_io_managers_0_grant_bits_is_builtin_type;
  wire [3:0] l1tol2net_io_managers_0_grant_bits_g_type;
  wire [63:0] l1tol2net_io_managers_0_grant_bits_data;
  wire  l1tol2net_io_managers_0_grant_bits_client_id;
  wire  l1tol2net_io_managers_0_finish_ready;
  wire  l1tol2net_io_managers_0_finish_valid;
  wire [1:0] l1tol2net_io_managers_0_finish_bits_manager_xact_id;
  wire  l1tol2net_io_managers_0_probe_ready;
  wire  l1tol2net_io_managers_0_probe_valid;
  wire [25:0] l1tol2net_io_managers_0_probe_bits_addr_block;
  wire [1:0] l1tol2net_io_managers_0_probe_bits_p_type;
  wire  l1tol2net_io_managers_0_probe_bits_client_id;
  wire  l1tol2net_io_managers_0_release_ready;
  wire  l1tol2net_io_managers_0_release_valid;
  wire [2:0] l1tol2net_io_managers_0_release_bits_addr_beat;
  wire [25:0] l1tol2net_io_managers_0_release_bits_addr_block;
  wire  l1tol2net_io_managers_0_release_bits_client_xact_id;
  wire  l1tol2net_io_managers_0_release_bits_voluntary;
  wire [2:0] l1tol2net_io_managers_0_release_bits_r_type;
  wire [63:0] l1tol2net_io_managers_0_release_bits_data;
  wire  l1tol2net_io_managers_0_release_bits_client_id;
  wire  l1tol2net_io_managers_1_acquire_ready;
  wire  l1tol2net_io_managers_1_acquire_valid;
  wire [25:0] l1tol2net_io_managers_1_acquire_bits_addr_block;
  wire  l1tol2net_io_managers_1_acquire_bits_client_xact_id;
  wire [2:0] l1tol2net_io_managers_1_acquire_bits_addr_beat;
  wire  l1tol2net_io_managers_1_acquire_bits_is_builtin_type;
  wire [2:0] l1tol2net_io_managers_1_acquire_bits_a_type;
  wire [11:0] l1tol2net_io_managers_1_acquire_bits_union;
  wire [63:0] l1tol2net_io_managers_1_acquire_bits_data;
  wire  l1tol2net_io_managers_1_acquire_bits_client_id;
  wire  l1tol2net_io_managers_1_grant_ready;
  wire  l1tol2net_io_managers_1_grant_valid;
  wire [2:0] l1tol2net_io_managers_1_grant_bits_addr_beat;
  wire  l1tol2net_io_managers_1_grant_bits_client_xact_id;
  wire [1:0] l1tol2net_io_managers_1_grant_bits_manager_xact_id;
  wire  l1tol2net_io_managers_1_grant_bits_is_builtin_type;
  wire [3:0] l1tol2net_io_managers_1_grant_bits_g_type;
  wire [63:0] l1tol2net_io_managers_1_grant_bits_data;
  wire  l1tol2net_io_managers_1_grant_bits_client_id;
  wire  l1tol2net_io_managers_1_finish_ready;
  wire  l1tol2net_io_managers_1_finish_valid;
  wire [1:0] l1tol2net_io_managers_1_finish_bits_manager_xact_id;
  wire  l1tol2net_io_managers_1_probe_ready;
  wire  l1tol2net_io_managers_1_probe_valid;
  wire [25:0] l1tol2net_io_managers_1_probe_bits_addr_block;
  wire [1:0] l1tol2net_io_managers_1_probe_bits_p_type;
  wire  l1tol2net_io_managers_1_probe_bits_client_id;
  wire  l1tol2net_io_managers_1_release_ready;
  wire  l1tol2net_io_managers_1_release_valid;
  wire [2:0] l1tol2net_io_managers_1_release_bits_addr_beat;
  wire [25:0] l1tol2net_io_managers_1_release_bits_addr_block;
  wire  l1tol2net_io_managers_1_release_bits_client_xact_id;
  wire  l1tol2net_io_managers_1_release_bits_voluntary;
  wire [2:0] l1tol2net_io_managers_1_release_bits_r_type;
  wire [63:0] l1tol2net_io_managers_1_release_bits_data;
  wire  l1tol2net_io_managers_1_release_bits_client_id;
  wire  ManagerToClientStatelessBridge_1_clk;
  wire  ManagerToClientStatelessBridge_1_reset;
  wire  ManagerToClientStatelessBridge_1_io_inner_acquire_ready;
  wire  ManagerToClientStatelessBridge_1_io_inner_acquire_valid;
  wire [25:0] ManagerToClientStatelessBridge_1_io_inner_acquire_bits_addr_block;
  wire  ManagerToClientStatelessBridge_1_io_inner_acquire_bits_client_xact_id;
  wire [2:0] ManagerToClientStatelessBridge_1_io_inner_acquire_bits_addr_beat;
  wire  ManagerToClientStatelessBridge_1_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] ManagerToClientStatelessBridge_1_io_inner_acquire_bits_a_type;
  wire [11:0] ManagerToClientStatelessBridge_1_io_inner_acquire_bits_union;
  wire [63:0] ManagerToClientStatelessBridge_1_io_inner_acquire_bits_data;
  wire  ManagerToClientStatelessBridge_1_io_inner_acquire_bits_client_id;
  wire  ManagerToClientStatelessBridge_1_io_inner_grant_ready;
  wire  ManagerToClientStatelessBridge_1_io_inner_grant_valid;
  wire [2:0] ManagerToClientStatelessBridge_1_io_inner_grant_bits_addr_beat;
  wire  ManagerToClientStatelessBridge_1_io_inner_grant_bits_client_xact_id;
  wire [1:0] ManagerToClientStatelessBridge_1_io_inner_grant_bits_manager_xact_id;
  wire  ManagerToClientStatelessBridge_1_io_inner_grant_bits_is_builtin_type;
  wire [3:0] ManagerToClientStatelessBridge_1_io_inner_grant_bits_g_type;
  wire [63:0] ManagerToClientStatelessBridge_1_io_inner_grant_bits_data;
  wire  ManagerToClientStatelessBridge_1_io_inner_grant_bits_client_id;
  wire  ManagerToClientStatelessBridge_1_io_inner_finish_ready;
  wire  ManagerToClientStatelessBridge_1_io_inner_finish_valid;
  wire [1:0] ManagerToClientStatelessBridge_1_io_inner_finish_bits_manager_xact_id;
  wire  ManagerToClientStatelessBridge_1_io_inner_probe_ready;
  wire  ManagerToClientStatelessBridge_1_io_inner_probe_valid;
  wire [25:0] ManagerToClientStatelessBridge_1_io_inner_probe_bits_addr_block;
  wire [1:0] ManagerToClientStatelessBridge_1_io_inner_probe_bits_p_type;
  wire  ManagerToClientStatelessBridge_1_io_inner_probe_bits_client_id;
  wire  ManagerToClientStatelessBridge_1_io_inner_release_ready;
  wire  ManagerToClientStatelessBridge_1_io_inner_release_valid;
  wire [2:0] ManagerToClientStatelessBridge_1_io_inner_release_bits_addr_beat;
  wire [25:0] ManagerToClientStatelessBridge_1_io_inner_release_bits_addr_block;
  wire  ManagerToClientStatelessBridge_1_io_inner_release_bits_client_xact_id;
  wire  ManagerToClientStatelessBridge_1_io_inner_release_bits_voluntary;
  wire [2:0] ManagerToClientStatelessBridge_1_io_inner_release_bits_r_type;
  wire [63:0] ManagerToClientStatelessBridge_1_io_inner_release_bits_data;
  wire  ManagerToClientStatelessBridge_1_io_inner_release_bits_client_id;
  wire  ManagerToClientStatelessBridge_1_io_incoherent_0;
  wire  ManagerToClientStatelessBridge_1_io_outer_acquire_ready;
  wire  ManagerToClientStatelessBridge_1_io_outer_acquire_valid;
  wire [25:0] ManagerToClientStatelessBridge_1_io_outer_acquire_bits_addr_block;
  wire [1:0] ManagerToClientStatelessBridge_1_io_outer_acquire_bits_client_xact_id;
  wire [2:0] ManagerToClientStatelessBridge_1_io_outer_acquire_bits_addr_beat;
  wire  ManagerToClientStatelessBridge_1_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] ManagerToClientStatelessBridge_1_io_outer_acquire_bits_a_type;
  wire [11:0] ManagerToClientStatelessBridge_1_io_outer_acquire_bits_union;
  wire [63:0] ManagerToClientStatelessBridge_1_io_outer_acquire_bits_data;
  wire  ManagerToClientStatelessBridge_1_io_outer_probe_ready;
  wire  ManagerToClientStatelessBridge_1_io_outer_probe_valid;
  wire [25:0] ManagerToClientStatelessBridge_1_io_outer_probe_bits_addr_block;
  wire [1:0] ManagerToClientStatelessBridge_1_io_outer_probe_bits_p_type;
  wire  ManagerToClientStatelessBridge_1_io_outer_release_ready;
  wire  ManagerToClientStatelessBridge_1_io_outer_release_valid;
  wire [2:0] ManagerToClientStatelessBridge_1_io_outer_release_bits_addr_beat;
  wire [25:0] ManagerToClientStatelessBridge_1_io_outer_release_bits_addr_block;
  wire [1:0] ManagerToClientStatelessBridge_1_io_outer_release_bits_client_xact_id;
  wire  ManagerToClientStatelessBridge_1_io_outer_release_bits_voluntary;
  wire [2:0] ManagerToClientStatelessBridge_1_io_outer_release_bits_r_type;
  wire [63:0] ManagerToClientStatelessBridge_1_io_outer_release_bits_data;
  wire  ManagerToClientStatelessBridge_1_io_outer_grant_ready;
  wire  ManagerToClientStatelessBridge_1_io_outer_grant_valid;
  wire [2:0] ManagerToClientStatelessBridge_1_io_outer_grant_bits_addr_beat;
  wire [1:0] ManagerToClientStatelessBridge_1_io_outer_grant_bits_client_xact_id;
  wire  ManagerToClientStatelessBridge_1_io_outer_grant_bits_manager_xact_id;
  wire  ManagerToClientStatelessBridge_1_io_outer_grant_bits_is_builtin_type;
  wire [3:0] ManagerToClientStatelessBridge_1_io_outer_grant_bits_g_type;
  wire [63:0] ManagerToClientStatelessBridge_1_io_outer_grant_bits_data;
  wire  ManagerToClientStatelessBridge_1_io_outer_grant_bits_manager_id;
  wire  ManagerToClientStatelessBridge_1_io_outer_finish_ready;
  wire  ManagerToClientStatelessBridge_1_io_outer_finish_valid;
  wire  ManagerToClientStatelessBridge_1_io_outer_finish_bits_manager_xact_id;
  wire  ManagerToClientStatelessBridge_1_io_outer_finish_bits_manager_id;
  wire  mmioManager_clk;
  wire  mmioManager_reset;
  wire  mmioManager_io_inner_acquire_ready;
  wire  mmioManager_io_inner_acquire_valid;
  wire [25:0] mmioManager_io_inner_acquire_bits_addr_block;
  wire  mmioManager_io_inner_acquire_bits_client_xact_id;
  wire [2:0] mmioManager_io_inner_acquire_bits_addr_beat;
  wire  mmioManager_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] mmioManager_io_inner_acquire_bits_a_type;
  wire [11:0] mmioManager_io_inner_acquire_bits_union;
  wire [63:0] mmioManager_io_inner_acquire_bits_data;
  wire  mmioManager_io_inner_acquire_bits_client_id;
  wire  mmioManager_io_inner_grant_ready;
  wire  mmioManager_io_inner_grant_valid;
  wire [2:0] mmioManager_io_inner_grant_bits_addr_beat;
  wire  mmioManager_io_inner_grant_bits_client_xact_id;
  wire [1:0] mmioManager_io_inner_grant_bits_manager_xact_id;
  wire  mmioManager_io_inner_grant_bits_is_builtin_type;
  wire [3:0] mmioManager_io_inner_grant_bits_g_type;
  wire [63:0] mmioManager_io_inner_grant_bits_data;
  wire  mmioManager_io_inner_grant_bits_client_id;
  wire  mmioManager_io_inner_finish_ready;
  wire  mmioManager_io_inner_finish_valid;
  wire [1:0] mmioManager_io_inner_finish_bits_manager_xact_id;
  wire  mmioManager_io_inner_probe_ready;
  wire  mmioManager_io_inner_probe_valid;
  wire [25:0] mmioManager_io_inner_probe_bits_addr_block;
  wire [1:0] mmioManager_io_inner_probe_bits_p_type;
  wire  mmioManager_io_inner_probe_bits_client_id;
  wire  mmioManager_io_inner_release_ready;
  wire  mmioManager_io_inner_release_valid;
  wire [2:0] mmioManager_io_inner_release_bits_addr_beat;
  wire [25:0] mmioManager_io_inner_release_bits_addr_block;
  wire  mmioManager_io_inner_release_bits_client_xact_id;
  wire  mmioManager_io_inner_release_bits_voluntary;
  wire [2:0] mmioManager_io_inner_release_bits_r_type;
  wire [63:0] mmioManager_io_inner_release_bits_data;
  wire  mmioManager_io_inner_release_bits_client_id;
  wire  mmioManager_io_incoherent_0;
  wire  mmioManager_io_outer_acquire_ready;
  wire  mmioManager_io_outer_acquire_valid;
  wire [25:0] mmioManager_io_outer_acquire_bits_addr_block;
  wire [1:0] mmioManager_io_outer_acquire_bits_client_xact_id;
  wire [2:0] mmioManager_io_outer_acquire_bits_addr_beat;
  wire  mmioManager_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] mmioManager_io_outer_acquire_bits_a_type;
  wire [11:0] mmioManager_io_outer_acquire_bits_union;
  wire [63:0] mmioManager_io_outer_acquire_bits_data;
  wire  mmioManager_io_outer_grant_ready;
  wire  mmioManager_io_outer_grant_valid;
  wire [2:0] mmioManager_io_outer_grant_bits_addr_beat;
  wire [1:0] mmioManager_io_outer_grant_bits_client_xact_id;
  wire  mmioManager_io_outer_grant_bits_manager_xact_id;
  wire  mmioManager_io_outer_grant_bits_is_builtin_type;
  wire [3:0] mmioManager_io_outer_grant_bits_g_type;
  wire [63:0] mmioManager_io_outer_grant_bits_data;
  wire  Queue_8_1_clk;
  wire  Queue_8_1_reset;
  wire  Queue_8_1_io_enq_ready;
  wire  Queue_8_1_io_enq_valid;
  wire [25:0] Queue_8_1_io_enq_bits_addr_block;
  wire [1:0] Queue_8_1_io_enq_bits_client_xact_id;
  wire [2:0] Queue_8_1_io_enq_bits_addr_beat;
  wire  Queue_8_1_io_enq_bits_is_builtin_type;
  wire [2:0] Queue_8_1_io_enq_bits_a_type;
  wire [11:0] Queue_8_1_io_enq_bits_union;
  wire [63:0] Queue_8_1_io_enq_bits_data;
  wire  Queue_8_1_io_deq_ready;
  wire  Queue_8_1_io_deq_valid;
  wire [25:0] Queue_8_1_io_deq_bits_addr_block;
  wire [1:0] Queue_8_1_io_deq_bits_client_xact_id;
  wire [2:0] Queue_8_1_io_deq_bits_addr_beat;
  wire  Queue_8_1_io_deq_bits_is_builtin_type;
  wire [2:0] Queue_8_1_io_deq_bits_a_type;
  wire [11:0] Queue_8_1_io_deq_bits_union;
  wire [63:0] Queue_8_1_io_deq_bits_data;
  wire  Queue_8_1_io_count;
  wire  Queue_9_1_clk;
  wire  Queue_9_1_reset;
  wire  Queue_9_1_io_enq_ready;
  wire  Queue_9_1_io_enq_valid;
  wire [2:0] Queue_9_1_io_enq_bits_addr_beat;
  wire [1:0] Queue_9_1_io_enq_bits_client_xact_id;
  wire  Queue_9_1_io_enq_bits_manager_xact_id;
  wire  Queue_9_1_io_enq_bits_is_builtin_type;
  wire [3:0] Queue_9_1_io_enq_bits_g_type;
  wire [63:0] Queue_9_1_io_enq_bits_data;
  wire  Queue_9_1_io_deq_ready;
  wire  Queue_9_1_io_deq_valid;
  wire [2:0] Queue_9_1_io_deq_bits_addr_beat;
  wire [1:0] Queue_9_1_io_deq_bits_client_xact_id;
  wire  Queue_9_1_io_deq_bits_manager_xact_id;
  wire  Queue_9_1_io_deq_bits_is_builtin_type;
  wire [3:0] Queue_9_1_io_deq_bits_g_type;
  wire [63:0] Queue_9_1_io_deq_bits_data;
  wire  Queue_9_1_io_count;
  wire  mem_ic_clk;
  wire  mem_ic_reset;
  wire  mem_ic_io_in_0_acquire_ready;
  wire  mem_ic_io_in_0_acquire_valid;
  wire [25:0] mem_ic_io_in_0_acquire_bits_addr_block;
  wire [1:0] mem_ic_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] mem_ic_io_in_0_acquire_bits_addr_beat;
  wire  mem_ic_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] mem_ic_io_in_0_acquire_bits_a_type;
  wire [11:0] mem_ic_io_in_0_acquire_bits_union;
  wire [63:0] mem_ic_io_in_0_acquire_bits_data;
  wire  mem_ic_io_in_0_grant_ready;
  wire  mem_ic_io_in_0_grant_valid;
  wire [2:0] mem_ic_io_in_0_grant_bits_addr_beat;
  wire [1:0] mem_ic_io_in_0_grant_bits_client_xact_id;
  wire  mem_ic_io_in_0_grant_bits_manager_xact_id;
  wire  mem_ic_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] mem_ic_io_in_0_grant_bits_g_type;
  wire [63:0] mem_ic_io_in_0_grant_bits_data;
  wire  mem_ic_io_out_0_acquire_ready;
  wire  mem_ic_io_out_0_acquire_valid;
  wire [25:0] mem_ic_io_out_0_acquire_bits_addr_block;
  wire [1:0] mem_ic_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] mem_ic_io_out_0_acquire_bits_addr_beat;
  wire  mem_ic_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] mem_ic_io_out_0_acquire_bits_a_type;
  wire [11:0] mem_ic_io_out_0_acquire_bits_union;
  wire [63:0] mem_ic_io_out_0_acquire_bits_data;
  wire  mem_ic_io_out_0_grant_ready;
  wire  mem_ic_io_out_0_grant_valid;
  wire [2:0] mem_ic_io_out_0_grant_bits_addr_beat;
  wire [1:0] mem_ic_io_out_0_grant_bits_client_xact_id;
  wire  mem_ic_io_out_0_grant_bits_manager_xact_id;
  wire  mem_ic_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] mem_ic_io_out_0_grant_bits_g_type;
  wire [63:0] mem_ic_io_out_0_grant_bits_data;
  wire  ClientTileLinkIOUnwrapper_1_clk;
  wire  ClientTileLinkIOUnwrapper_1_reset;
  wire  ClientTileLinkIOUnwrapper_1_io_in_acquire_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_in_acquire_valid;
  wire [25:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_block;
  wire [1:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_beat;
  wire  ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_a_type;
  wire [11:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_union;
  wire [63:0] ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_data;
  wire  ClientTileLinkIOUnwrapper_1_io_in_probe_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_in_probe_valid;
  wire [25:0] ClientTileLinkIOUnwrapper_1_io_in_probe_bits_addr_block;
  wire [1:0] ClientTileLinkIOUnwrapper_1_io_in_probe_bits_p_type;
  wire  ClientTileLinkIOUnwrapper_1_io_in_release_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_in_release_valid;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_beat;
  wire [25:0] ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_block;
  wire [1:0] ClientTileLinkIOUnwrapper_1_io_in_release_bits_client_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_in_release_bits_voluntary;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_release_bits_r_type;
  wire [63:0] ClientTileLinkIOUnwrapper_1_io_in_release_bits_data;
  wire  ClientTileLinkIOUnwrapper_1_io_in_grant_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_in_grant_valid;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_in_grant_bits_addr_beat;
  wire [1:0] ClientTileLinkIOUnwrapper_1_io_in_grant_bits_client_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_in_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkIOUnwrapper_1_io_in_grant_bits_g_type;
  wire [63:0] ClientTileLinkIOUnwrapper_1_io_in_grant_bits_data;
  wire  ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_id;
  wire  ClientTileLinkIOUnwrapper_1_io_in_finish_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_in_finish_valid;
  wire  ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_id;
  wire  ClientTileLinkIOUnwrapper_1_io_out_acquire_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_out_acquire_valid;
  wire [25:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_block;
  wire [1:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_beat;
  wire  ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_a_type;
  wire [11:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_union;
  wire [63:0] ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_data;
  wire  ClientTileLinkIOUnwrapper_1_io_out_grant_ready;
  wire  ClientTileLinkIOUnwrapper_1_io_out_grant_valid;
  wire [2:0] ClientTileLinkIOUnwrapper_1_io_out_grant_bits_addr_beat;
  wire [1:0] ClientTileLinkIOUnwrapper_1_io_out_grant_bits_client_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_out_grant_bits_manager_xact_id;
  wire  ClientTileLinkIOUnwrapper_1_io_out_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkIOUnwrapper_1_io_out_grant_bits_g_type;
  wire [63:0] ClientTileLinkIOUnwrapper_1_io_out_grant_bits_data;
  wire  ClientTileLinkEnqueuer_1_clk;
  wire  ClientTileLinkEnqueuer_1_reset;
  wire  ClientTileLinkEnqueuer_1_io_inner_acquire_ready;
  wire  ClientTileLinkEnqueuer_1_io_inner_acquire_valid;
  wire [25:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_block;
  wire [1:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_beat;
  wire  ClientTileLinkEnqueuer_1_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_a_type;
  wire [11:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_union;
  wire [63:0] ClientTileLinkEnqueuer_1_io_inner_acquire_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_inner_probe_ready;
  wire  ClientTileLinkEnqueuer_1_io_inner_probe_valid;
  wire [25:0] ClientTileLinkEnqueuer_1_io_inner_probe_bits_addr_block;
  wire [1:0] ClientTileLinkEnqueuer_1_io_inner_probe_bits_p_type;
  wire  ClientTileLinkEnqueuer_1_io_inner_release_ready;
  wire  ClientTileLinkEnqueuer_1_io_inner_release_valid;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_beat;
  wire [25:0] ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_block;
  wire [1:0] ClientTileLinkEnqueuer_1_io_inner_release_bits_client_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_inner_release_bits_voluntary;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_release_bits_r_type;
  wire [63:0] ClientTileLinkEnqueuer_1_io_inner_release_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_inner_grant_ready;
  wire  ClientTileLinkEnqueuer_1_io_inner_grant_valid;
  wire [2:0] ClientTileLinkEnqueuer_1_io_inner_grant_bits_addr_beat;
  wire [1:0] ClientTileLinkEnqueuer_1_io_inner_grant_bits_client_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_inner_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkEnqueuer_1_io_inner_grant_bits_g_type;
  wire [63:0] ClientTileLinkEnqueuer_1_io_inner_grant_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_id;
  wire  ClientTileLinkEnqueuer_1_io_inner_finish_ready;
  wire  ClientTileLinkEnqueuer_1_io_inner_finish_valid;
  wire  ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_acquire_ready;
  wire  ClientTileLinkEnqueuer_1_io_outer_acquire_valid;
  wire [25:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_block;
  wire [1:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_beat;
  wire  ClientTileLinkEnqueuer_1_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_a_type;
  wire [11:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_union;
  wire [63:0] ClientTileLinkEnqueuer_1_io_outer_acquire_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_outer_probe_ready;
  wire  ClientTileLinkEnqueuer_1_io_outer_probe_valid;
  wire [25:0] ClientTileLinkEnqueuer_1_io_outer_probe_bits_addr_block;
  wire [1:0] ClientTileLinkEnqueuer_1_io_outer_probe_bits_p_type;
  wire  ClientTileLinkEnqueuer_1_io_outer_release_ready;
  wire  ClientTileLinkEnqueuer_1_io_outer_release_valid;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_beat;
  wire [25:0] ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_block;
  wire [1:0] ClientTileLinkEnqueuer_1_io_outer_release_bits_client_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_release_bits_voluntary;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_release_bits_r_type;
  wire [63:0] ClientTileLinkEnqueuer_1_io_outer_release_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_outer_grant_ready;
  wire  ClientTileLinkEnqueuer_1_io_outer_grant_valid;
  wire [2:0] ClientTileLinkEnqueuer_1_io_outer_grant_bits_addr_beat;
  wire [1:0] ClientTileLinkEnqueuer_1_io_outer_grant_bits_client_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkEnqueuer_1_io_outer_grant_bits_g_type;
  wire [63:0] ClientTileLinkEnqueuer_1_io_outer_grant_bits_data;
  wire  ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_finish_ready;
  wire  ClientTileLinkEnqueuer_1_io_outer_finish_valid;
  wire  ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_xact_id;
  wire  ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_id;
  wire  NastiIOTileLinkIOConverter_1_clk;
  wire  NastiIOTileLinkIOConverter_1_reset;
  wire  NastiIOTileLinkIOConverter_1_io_tl_acquire_ready;
  wire  NastiIOTileLinkIOConverter_1_io_tl_acquire_valid;
  wire [25:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_block;
  wire [1:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_client_xact_id;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_beat;
  wire  NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_a_type;
  wire [11:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_union;
  wire [63:0] NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_data;
  wire  NastiIOTileLinkIOConverter_1_io_tl_grant_ready;
  wire  NastiIOTileLinkIOConverter_1_io_tl_grant_valid;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_tl_grant_bits_addr_beat;
  wire [1:0] NastiIOTileLinkIOConverter_1_io_tl_grant_bits_client_xact_id;
  wire  NastiIOTileLinkIOConverter_1_io_tl_grant_bits_manager_xact_id;
  wire  NastiIOTileLinkIOConverter_1_io_tl_grant_bits_is_builtin_type;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_tl_grant_bits_g_type;
  wire [63:0] NastiIOTileLinkIOConverter_1_io_tl_grant_bits_data;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_aw_ready;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_aw_valid;
  wire [31:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_addr;
  wire [7:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_len;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_size;
  wire [1:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_burst;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_lock;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_cache;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_prot;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_qos;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_region;
  wire [4:0] NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_id;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_user;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_w_ready;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_w_valid;
  wire [63:0] NastiIOTileLinkIOConverter_1_io_nasti_w_bits_data;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_w_bits_last;
  wire [4:0] NastiIOTileLinkIOConverter_1_io_nasti_w_bits_id;
  wire [7:0] NastiIOTileLinkIOConverter_1_io_nasti_w_bits_strb;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_w_bits_user;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_b_ready;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_b_valid;
  wire [1:0] NastiIOTileLinkIOConverter_1_io_nasti_b_bits_resp;
  wire [4:0] NastiIOTileLinkIOConverter_1_io_nasti_b_bits_id;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_b_bits_user;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_ar_ready;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_ar_valid;
  wire [31:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_addr;
  wire [7:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_len;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_size;
  wire [1:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_burst;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_lock;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_cache;
  wire [2:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_prot;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_qos;
  wire [3:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_region;
  wire [4:0] NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_id;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_user;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_r_ready;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_r_valid;
  wire [1:0] NastiIOTileLinkIOConverter_1_io_nasti_r_bits_resp;
  wire [63:0] NastiIOTileLinkIOConverter_1_io_nasti_r_bits_data;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_r_bits_last;
  wire [4:0] NastiIOTileLinkIOConverter_1_io_nasti_r_bits_id;
  wire  NastiIOTileLinkIOConverter_1_io_nasti_r_bits_user;
  wire  Queue_10_1_clk;
  wire  Queue_10_1_reset;
  wire  Queue_10_1_io_enq_ready;
  wire  Queue_10_1_io_enq_valid;
  wire [31:0] Queue_10_1_io_enq_bits_addr;
  wire [7:0] Queue_10_1_io_enq_bits_len;
  wire [2:0] Queue_10_1_io_enq_bits_size;
  wire [1:0] Queue_10_1_io_enq_bits_burst;
  wire  Queue_10_1_io_enq_bits_lock;
  wire [3:0] Queue_10_1_io_enq_bits_cache;
  wire [2:0] Queue_10_1_io_enq_bits_prot;
  wire [3:0] Queue_10_1_io_enq_bits_qos;
  wire [3:0] Queue_10_1_io_enq_bits_region;
  wire [4:0] Queue_10_1_io_enq_bits_id;
  wire  Queue_10_1_io_enq_bits_user;
  wire  Queue_10_1_io_deq_ready;
  wire  Queue_10_1_io_deq_valid;
  wire [31:0] Queue_10_1_io_deq_bits_addr;
  wire [7:0] Queue_10_1_io_deq_bits_len;
  wire [2:0] Queue_10_1_io_deq_bits_size;
  wire [1:0] Queue_10_1_io_deq_bits_burst;
  wire  Queue_10_1_io_deq_bits_lock;
  wire [3:0] Queue_10_1_io_deq_bits_cache;
  wire [2:0] Queue_10_1_io_deq_bits_prot;
  wire [3:0] Queue_10_1_io_deq_bits_qos;
  wire [3:0] Queue_10_1_io_deq_bits_region;
  wire [4:0] Queue_10_1_io_deq_bits_id;
  wire  Queue_10_1_io_deq_bits_user;
  wire  Queue_10_1_io_count;
  wire  Queue_11_1_clk;
  wire  Queue_11_1_reset;
  wire  Queue_11_1_io_enq_ready;
  wire  Queue_11_1_io_enq_valid;
  wire [31:0] Queue_11_1_io_enq_bits_addr;
  wire [7:0] Queue_11_1_io_enq_bits_len;
  wire [2:0] Queue_11_1_io_enq_bits_size;
  wire [1:0] Queue_11_1_io_enq_bits_burst;
  wire  Queue_11_1_io_enq_bits_lock;
  wire [3:0] Queue_11_1_io_enq_bits_cache;
  wire [2:0] Queue_11_1_io_enq_bits_prot;
  wire [3:0] Queue_11_1_io_enq_bits_qos;
  wire [3:0] Queue_11_1_io_enq_bits_region;
  wire [4:0] Queue_11_1_io_enq_bits_id;
  wire  Queue_11_1_io_enq_bits_user;
  wire  Queue_11_1_io_deq_ready;
  wire  Queue_11_1_io_deq_valid;
  wire [31:0] Queue_11_1_io_deq_bits_addr;
  wire [7:0] Queue_11_1_io_deq_bits_len;
  wire [2:0] Queue_11_1_io_deq_bits_size;
  wire [1:0] Queue_11_1_io_deq_bits_burst;
  wire  Queue_11_1_io_deq_bits_lock;
  wire [3:0] Queue_11_1_io_deq_bits_cache;
  wire [2:0] Queue_11_1_io_deq_bits_prot;
  wire [3:0] Queue_11_1_io_deq_bits_qos;
  wire [3:0] Queue_11_1_io_deq_bits_region;
  wire [4:0] Queue_11_1_io_deq_bits_id;
  wire  Queue_11_1_io_deq_bits_user;
  wire  Queue_11_1_io_count;
  wire  Queue_12_1_clk;
  wire  Queue_12_1_reset;
  wire  Queue_12_1_io_enq_ready;
  wire  Queue_12_1_io_enq_valid;
  wire [63:0] Queue_12_1_io_enq_bits_data;
  wire  Queue_12_1_io_enq_bits_last;
  wire [4:0] Queue_12_1_io_enq_bits_id;
  wire [7:0] Queue_12_1_io_enq_bits_strb;
  wire  Queue_12_1_io_enq_bits_user;
  wire  Queue_12_1_io_deq_ready;
  wire  Queue_12_1_io_deq_valid;
  wire [63:0] Queue_12_1_io_deq_bits_data;
  wire  Queue_12_1_io_deq_bits_last;
  wire [4:0] Queue_12_1_io_deq_bits_id;
  wire [7:0] Queue_12_1_io_deq_bits_strb;
  wire  Queue_12_1_io_deq_bits_user;
  wire [1:0] Queue_12_1_io_count;
  wire  Queue_13_1_clk;
  wire  Queue_13_1_reset;
  wire  Queue_13_1_io_enq_ready;
  wire  Queue_13_1_io_enq_valid;
  wire [1:0] Queue_13_1_io_enq_bits_resp;
  wire [63:0] Queue_13_1_io_enq_bits_data;
  wire  Queue_13_1_io_enq_bits_last;
  wire [4:0] Queue_13_1_io_enq_bits_id;
  wire  Queue_13_1_io_enq_bits_user;
  wire  Queue_13_1_io_deq_ready;
  wire  Queue_13_1_io_deq_valid;
  wire [1:0] Queue_13_1_io_deq_bits_resp;
  wire [63:0] Queue_13_1_io_deq_bits_data;
  wire  Queue_13_1_io_deq_bits_last;
  wire [4:0] Queue_13_1_io_deq_bits_id;
  wire  Queue_13_1_io_deq_bits_user;
  wire [1:0] Queue_13_1_io_count;
  wire  Queue_14_1_clk;
  wire  Queue_14_1_reset;
  wire  Queue_14_1_io_enq_ready;
  wire  Queue_14_1_io_enq_valid;
  wire [1:0] Queue_14_1_io_enq_bits_resp;
  wire [4:0] Queue_14_1_io_enq_bits_id;
  wire  Queue_14_1_io_enq_bits_user;
  wire  Queue_14_1_io_deq_ready;
  wire  Queue_14_1_io_deq_valid;
  wire [1:0] Queue_14_1_io_deq_bits_resp;
  wire [4:0] Queue_14_1_io_deq_bits_id;
  wire  Queue_14_1_io_deq_bits_user;
  wire  Queue_14_1_io_count;
  reg  GEN_0;
  reg [31:0] GEN_1;
  PortedTileLinkCrossbar l1tol2net (
    .clk(l1tol2net_clk),
    .reset(l1tol2net_reset),
    .io_clients_cached_0_acquire_ready(l1tol2net_io_clients_cached_0_acquire_ready),
    .io_clients_cached_0_acquire_valid(l1tol2net_io_clients_cached_0_acquire_valid),
    .io_clients_cached_0_acquire_bits_addr_block(l1tol2net_io_clients_cached_0_acquire_bits_addr_block),
    .io_clients_cached_0_acquire_bits_client_xact_id(l1tol2net_io_clients_cached_0_acquire_bits_client_xact_id),
    .io_clients_cached_0_acquire_bits_addr_beat(l1tol2net_io_clients_cached_0_acquire_bits_addr_beat),
    .io_clients_cached_0_acquire_bits_is_builtin_type(l1tol2net_io_clients_cached_0_acquire_bits_is_builtin_type),
    .io_clients_cached_0_acquire_bits_a_type(l1tol2net_io_clients_cached_0_acquire_bits_a_type),
    .io_clients_cached_0_acquire_bits_union(l1tol2net_io_clients_cached_0_acquire_bits_union),
    .io_clients_cached_0_acquire_bits_data(l1tol2net_io_clients_cached_0_acquire_bits_data),
    .io_clients_cached_0_probe_ready(l1tol2net_io_clients_cached_0_probe_ready),
    .io_clients_cached_0_probe_valid(l1tol2net_io_clients_cached_0_probe_valid),
    .io_clients_cached_0_probe_bits_addr_block(l1tol2net_io_clients_cached_0_probe_bits_addr_block),
    .io_clients_cached_0_probe_bits_p_type(l1tol2net_io_clients_cached_0_probe_bits_p_type),
    .io_clients_cached_0_release_ready(l1tol2net_io_clients_cached_0_release_ready),
    .io_clients_cached_0_release_valid(l1tol2net_io_clients_cached_0_release_valid),
    .io_clients_cached_0_release_bits_addr_beat(l1tol2net_io_clients_cached_0_release_bits_addr_beat),
    .io_clients_cached_0_release_bits_addr_block(l1tol2net_io_clients_cached_0_release_bits_addr_block),
    .io_clients_cached_0_release_bits_client_xact_id(l1tol2net_io_clients_cached_0_release_bits_client_xact_id),
    .io_clients_cached_0_release_bits_voluntary(l1tol2net_io_clients_cached_0_release_bits_voluntary),
    .io_clients_cached_0_release_bits_r_type(l1tol2net_io_clients_cached_0_release_bits_r_type),
    .io_clients_cached_0_release_bits_data(l1tol2net_io_clients_cached_0_release_bits_data),
    .io_clients_cached_0_grant_ready(l1tol2net_io_clients_cached_0_grant_ready),
    .io_clients_cached_0_grant_valid(l1tol2net_io_clients_cached_0_grant_valid),
    .io_clients_cached_0_grant_bits_addr_beat(l1tol2net_io_clients_cached_0_grant_bits_addr_beat),
    .io_clients_cached_0_grant_bits_client_xact_id(l1tol2net_io_clients_cached_0_grant_bits_client_xact_id),
    .io_clients_cached_0_grant_bits_manager_xact_id(l1tol2net_io_clients_cached_0_grant_bits_manager_xact_id),
    .io_clients_cached_0_grant_bits_is_builtin_type(l1tol2net_io_clients_cached_0_grant_bits_is_builtin_type),
    .io_clients_cached_0_grant_bits_g_type(l1tol2net_io_clients_cached_0_grant_bits_g_type),
    .io_clients_cached_0_grant_bits_data(l1tol2net_io_clients_cached_0_grant_bits_data),
    .io_clients_cached_0_grant_bits_manager_id(l1tol2net_io_clients_cached_0_grant_bits_manager_id),
    .io_clients_cached_0_finish_ready(l1tol2net_io_clients_cached_0_finish_ready),
    .io_clients_cached_0_finish_valid(l1tol2net_io_clients_cached_0_finish_valid),
    .io_clients_cached_0_finish_bits_manager_xact_id(l1tol2net_io_clients_cached_0_finish_bits_manager_xact_id),
    .io_clients_cached_0_finish_bits_manager_id(l1tol2net_io_clients_cached_0_finish_bits_manager_id),
    .io_clients_uncached_0_acquire_ready(l1tol2net_io_clients_uncached_0_acquire_ready),
    .io_clients_uncached_0_acquire_valid(l1tol2net_io_clients_uncached_0_acquire_valid),
    .io_clients_uncached_0_acquire_bits_addr_block(l1tol2net_io_clients_uncached_0_acquire_bits_addr_block),
    .io_clients_uncached_0_acquire_bits_client_xact_id(l1tol2net_io_clients_uncached_0_acquire_bits_client_xact_id),
    .io_clients_uncached_0_acquire_bits_addr_beat(l1tol2net_io_clients_uncached_0_acquire_bits_addr_beat),
    .io_clients_uncached_0_acquire_bits_is_builtin_type(l1tol2net_io_clients_uncached_0_acquire_bits_is_builtin_type),
    .io_clients_uncached_0_acquire_bits_a_type(l1tol2net_io_clients_uncached_0_acquire_bits_a_type),
    .io_clients_uncached_0_acquire_bits_union(l1tol2net_io_clients_uncached_0_acquire_bits_union),
    .io_clients_uncached_0_acquire_bits_data(l1tol2net_io_clients_uncached_0_acquire_bits_data),
    .io_clients_uncached_0_grant_ready(l1tol2net_io_clients_uncached_0_grant_ready),
    .io_clients_uncached_0_grant_valid(l1tol2net_io_clients_uncached_0_grant_valid),
    .io_clients_uncached_0_grant_bits_addr_beat(l1tol2net_io_clients_uncached_0_grant_bits_addr_beat),
    .io_clients_uncached_0_grant_bits_client_xact_id(l1tol2net_io_clients_uncached_0_grant_bits_client_xact_id),
    .io_clients_uncached_0_grant_bits_manager_xact_id(l1tol2net_io_clients_uncached_0_grant_bits_manager_xact_id),
    .io_clients_uncached_0_grant_bits_is_builtin_type(l1tol2net_io_clients_uncached_0_grant_bits_is_builtin_type),
    .io_clients_uncached_0_grant_bits_g_type(l1tol2net_io_clients_uncached_0_grant_bits_g_type),
    .io_clients_uncached_0_grant_bits_data(l1tol2net_io_clients_uncached_0_grant_bits_data),
    .io_managers_0_acquire_ready(l1tol2net_io_managers_0_acquire_ready),
    .io_managers_0_acquire_valid(l1tol2net_io_managers_0_acquire_valid),
    .io_managers_0_acquire_bits_addr_block(l1tol2net_io_managers_0_acquire_bits_addr_block),
    .io_managers_0_acquire_bits_client_xact_id(l1tol2net_io_managers_0_acquire_bits_client_xact_id),
    .io_managers_0_acquire_bits_addr_beat(l1tol2net_io_managers_0_acquire_bits_addr_beat),
    .io_managers_0_acquire_bits_is_builtin_type(l1tol2net_io_managers_0_acquire_bits_is_builtin_type),
    .io_managers_0_acquire_bits_a_type(l1tol2net_io_managers_0_acquire_bits_a_type),
    .io_managers_0_acquire_bits_union(l1tol2net_io_managers_0_acquire_bits_union),
    .io_managers_0_acquire_bits_data(l1tol2net_io_managers_0_acquire_bits_data),
    .io_managers_0_acquire_bits_client_id(l1tol2net_io_managers_0_acquire_bits_client_id),
    .io_managers_0_grant_ready(l1tol2net_io_managers_0_grant_ready),
    .io_managers_0_grant_valid(l1tol2net_io_managers_0_grant_valid),
    .io_managers_0_grant_bits_addr_beat(l1tol2net_io_managers_0_grant_bits_addr_beat),
    .io_managers_0_grant_bits_client_xact_id(l1tol2net_io_managers_0_grant_bits_client_xact_id),
    .io_managers_0_grant_bits_manager_xact_id(l1tol2net_io_managers_0_grant_bits_manager_xact_id),
    .io_managers_0_grant_bits_is_builtin_type(l1tol2net_io_managers_0_grant_bits_is_builtin_type),
    .io_managers_0_grant_bits_g_type(l1tol2net_io_managers_0_grant_bits_g_type),
    .io_managers_0_grant_bits_data(l1tol2net_io_managers_0_grant_bits_data),
    .io_managers_0_grant_bits_client_id(l1tol2net_io_managers_0_grant_bits_client_id),
    .io_managers_0_finish_ready(l1tol2net_io_managers_0_finish_ready),
    .io_managers_0_finish_valid(l1tol2net_io_managers_0_finish_valid),
    .io_managers_0_finish_bits_manager_xact_id(l1tol2net_io_managers_0_finish_bits_manager_xact_id),
    .io_managers_0_probe_ready(l1tol2net_io_managers_0_probe_ready),
    .io_managers_0_probe_valid(l1tol2net_io_managers_0_probe_valid),
    .io_managers_0_probe_bits_addr_block(l1tol2net_io_managers_0_probe_bits_addr_block),
    .io_managers_0_probe_bits_p_type(l1tol2net_io_managers_0_probe_bits_p_type),
    .io_managers_0_probe_bits_client_id(l1tol2net_io_managers_0_probe_bits_client_id),
    .io_managers_0_release_ready(l1tol2net_io_managers_0_release_ready),
    .io_managers_0_release_valid(l1tol2net_io_managers_0_release_valid),
    .io_managers_0_release_bits_addr_beat(l1tol2net_io_managers_0_release_bits_addr_beat),
    .io_managers_0_release_bits_addr_block(l1tol2net_io_managers_0_release_bits_addr_block),
    .io_managers_0_release_bits_client_xact_id(l1tol2net_io_managers_0_release_bits_client_xact_id),
    .io_managers_0_release_bits_voluntary(l1tol2net_io_managers_0_release_bits_voluntary),
    .io_managers_0_release_bits_r_type(l1tol2net_io_managers_0_release_bits_r_type),
    .io_managers_0_release_bits_data(l1tol2net_io_managers_0_release_bits_data),
    .io_managers_0_release_bits_client_id(l1tol2net_io_managers_0_release_bits_client_id),
    .io_managers_1_acquire_ready(l1tol2net_io_managers_1_acquire_ready),
    .io_managers_1_acquire_valid(l1tol2net_io_managers_1_acquire_valid),
    .io_managers_1_acquire_bits_addr_block(l1tol2net_io_managers_1_acquire_bits_addr_block),
    .io_managers_1_acquire_bits_client_xact_id(l1tol2net_io_managers_1_acquire_bits_client_xact_id),
    .io_managers_1_acquire_bits_addr_beat(l1tol2net_io_managers_1_acquire_bits_addr_beat),
    .io_managers_1_acquire_bits_is_builtin_type(l1tol2net_io_managers_1_acquire_bits_is_builtin_type),
    .io_managers_1_acquire_bits_a_type(l1tol2net_io_managers_1_acquire_bits_a_type),
    .io_managers_1_acquire_bits_union(l1tol2net_io_managers_1_acquire_bits_union),
    .io_managers_1_acquire_bits_data(l1tol2net_io_managers_1_acquire_bits_data),
    .io_managers_1_acquire_bits_client_id(l1tol2net_io_managers_1_acquire_bits_client_id),
    .io_managers_1_grant_ready(l1tol2net_io_managers_1_grant_ready),
    .io_managers_1_grant_valid(l1tol2net_io_managers_1_grant_valid),
    .io_managers_1_grant_bits_addr_beat(l1tol2net_io_managers_1_grant_bits_addr_beat),
    .io_managers_1_grant_bits_client_xact_id(l1tol2net_io_managers_1_grant_bits_client_xact_id),
    .io_managers_1_grant_bits_manager_xact_id(l1tol2net_io_managers_1_grant_bits_manager_xact_id),
    .io_managers_1_grant_bits_is_builtin_type(l1tol2net_io_managers_1_grant_bits_is_builtin_type),
    .io_managers_1_grant_bits_g_type(l1tol2net_io_managers_1_grant_bits_g_type),
    .io_managers_1_grant_bits_data(l1tol2net_io_managers_1_grant_bits_data),
    .io_managers_1_grant_bits_client_id(l1tol2net_io_managers_1_grant_bits_client_id),
    .io_managers_1_finish_ready(l1tol2net_io_managers_1_finish_ready),
    .io_managers_1_finish_valid(l1tol2net_io_managers_1_finish_valid),
    .io_managers_1_finish_bits_manager_xact_id(l1tol2net_io_managers_1_finish_bits_manager_xact_id),
    .io_managers_1_probe_ready(l1tol2net_io_managers_1_probe_ready),
    .io_managers_1_probe_valid(l1tol2net_io_managers_1_probe_valid),
    .io_managers_1_probe_bits_addr_block(l1tol2net_io_managers_1_probe_bits_addr_block),
    .io_managers_1_probe_bits_p_type(l1tol2net_io_managers_1_probe_bits_p_type),
    .io_managers_1_probe_bits_client_id(l1tol2net_io_managers_1_probe_bits_client_id),
    .io_managers_1_release_ready(l1tol2net_io_managers_1_release_ready),
    .io_managers_1_release_valid(l1tol2net_io_managers_1_release_valid),
    .io_managers_1_release_bits_addr_beat(l1tol2net_io_managers_1_release_bits_addr_beat),
    .io_managers_1_release_bits_addr_block(l1tol2net_io_managers_1_release_bits_addr_block),
    .io_managers_1_release_bits_client_xact_id(l1tol2net_io_managers_1_release_bits_client_xact_id),
    .io_managers_1_release_bits_voluntary(l1tol2net_io_managers_1_release_bits_voluntary),
    .io_managers_1_release_bits_r_type(l1tol2net_io_managers_1_release_bits_r_type),
    .io_managers_1_release_bits_data(l1tol2net_io_managers_1_release_bits_data),
    .io_managers_1_release_bits_client_id(l1tol2net_io_managers_1_release_bits_client_id)
  );
  ManagerToClientStatelessBridge ManagerToClientStatelessBridge_1 (
    .clk(ManagerToClientStatelessBridge_1_clk),
    .reset(ManagerToClientStatelessBridge_1_reset),
    .io_inner_acquire_ready(ManagerToClientStatelessBridge_1_io_inner_acquire_ready),
    .io_inner_acquire_valid(ManagerToClientStatelessBridge_1_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(ManagerToClientStatelessBridge_1_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(ManagerToClientStatelessBridge_1_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(ManagerToClientStatelessBridge_1_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(ManagerToClientStatelessBridge_1_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(ManagerToClientStatelessBridge_1_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(ManagerToClientStatelessBridge_1_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(ManagerToClientStatelessBridge_1_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(ManagerToClientStatelessBridge_1_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(ManagerToClientStatelessBridge_1_io_inner_grant_ready),
    .io_inner_grant_valid(ManagerToClientStatelessBridge_1_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(ManagerToClientStatelessBridge_1_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(ManagerToClientStatelessBridge_1_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(ManagerToClientStatelessBridge_1_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(ManagerToClientStatelessBridge_1_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(ManagerToClientStatelessBridge_1_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(ManagerToClientStatelessBridge_1_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(ManagerToClientStatelessBridge_1_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(ManagerToClientStatelessBridge_1_io_inner_finish_ready),
    .io_inner_finish_valid(ManagerToClientStatelessBridge_1_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(ManagerToClientStatelessBridge_1_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(ManagerToClientStatelessBridge_1_io_inner_probe_ready),
    .io_inner_probe_valid(ManagerToClientStatelessBridge_1_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(ManagerToClientStatelessBridge_1_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(ManagerToClientStatelessBridge_1_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(ManagerToClientStatelessBridge_1_io_inner_probe_bits_client_id),
    .io_inner_release_ready(ManagerToClientStatelessBridge_1_io_inner_release_ready),
    .io_inner_release_valid(ManagerToClientStatelessBridge_1_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(ManagerToClientStatelessBridge_1_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(ManagerToClientStatelessBridge_1_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(ManagerToClientStatelessBridge_1_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(ManagerToClientStatelessBridge_1_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(ManagerToClientStatelessBridge_1_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(ManagerToClientStatelessBridge_1_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(ManagerToClientStatelessBridge_1_io_inner_release_bits_client_id),
    .io_incoherent_0(ManagerToClientStatelessBridge_1_io_incoherent_0),
    .io_outer_acquire_ready(ManagerToClientStatelessBridge_1_io_outer_acquire_ready),
    .io_outer_acquire_valid(ManagerToClientStatelessBridge_1_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(ManagerToClientStatelessBridge_1_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(ManagerToClientStatelessBridge_1_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(ManagerToClientStatelessBridge_1_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(ManagerToClientStatelessBridge_1_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(ManagerToClientStatelessBridge_1_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(ManagerToClientStatelessBridge_1_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(ManagerToClientStatelessBridge_1_io_outer_acquire_bits_data),
    .io_outer_probe_ready(ManagerToClientStatelessBridge_1_io_outer_probe_ready),
    .io_outer_probe_valid(ManagerToClientStatelessBridge_1_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(ManagerToClientStatelessBridge_1_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(ManagerToClientStatelessBridge_1_io_outer_probe_bits_p_type),
    .io_outer_release_ready(ManagerToClientStatelessBridge_1_io_outer_release_ready),
    .io_outer_release_valid(ManagerToClientStatelessBridge_1_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(ManagerToClientStatelessBridge_1_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(ManagerToClientStatelessBridge_1_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(ManagerToClientStatelessBridge_1_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(ManagerToClientStatelessBridge_1_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(ManagerToClientStatelessBridge_1_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(ManagerToClientStatelessBridge_1_io_outer_release_bits_data),
    .io_outer_grant_ready(ManagerToClientStatelessBridge_1_io_outer_grant_ready),
    .io_outer_grant_valid(ManagerToClientStatelessBridge_1_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(ManagerToClientStatelessBridge_1_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(ManagerToClientStatelessBridge_1_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(ManagerToClientStatelessBridge_1_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(ManagerToClientStatelessBridge_1_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(ManagerToClientStatelessBridge_1_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(ManagerToClientStatelessBridge_1_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(ManagerToClientStatelessBridge_1_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(ManagerToClientStatelessBridge_1_io_outer_finish_ready),
    .io_outer_finish_valid(ManagerToClientStatelessBridge_1_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(ManagerToClientStatelessBridge_1_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(ManagerToClientStatelessBridge_1_io_outer_finish_bits_manager_id)
  );
  MMIOTileLinkManager mmioManager (
    .clk(mmioManager_clk),
    .reset(mmioManager_reset),
    .io_inner_acquire_ready(mmioManager_io_inner_acquire_ready),
    .io_inner_acquire_valid(mmioManager_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(mmioManager_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(mmioManager_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(mmioManager_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(mmioManager_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(mmioManager_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(mmioManager_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(mmioManager_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(mmioManager_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(mmioManager_io_inner_grant_ready),
    .io_inner_grant_valid(mmioManager_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(mmioManager_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(mmioManager_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(mmioManager_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(mmioManager_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(mmioManager_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(mmioManager_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(mmioManager_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(mmioManager_io_inner_finish_ready),
    .io_inner_finish_valid(mmioManager_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(mmioManager_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(mmioManager_io_inner_probe_ready),
    .io_inner_probe_valid(mmioManager_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(mmioManager_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(mmioManager_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(mmioManager_io_inner_probe_bits_client_id),
    .io_inner_release_ready(mmioManager_io_inner_release_ready),
    .io_inner_release_valid(mmioManager_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(mmioManager_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(mmioManager_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(mmioManager_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(mmioManager_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(mmioManager_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(mmioManager_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(mmioManager_io_inner_release_bits_client_id),
    .io_incoherent_0(mmioManager_io_incoherent_0),
    .io_outer_acquire_ready(mmioManager_io_outer_acquire_ready),
    .io_outer_acquire_valid(mmioManager_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(mmioManager_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(mmioManager_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(mmioManager_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(mmioManager_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(mmioManager_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(mmioManager_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(mmioManager_io_outer_acquire_bits_data),
    .io_outer_grant_ready(mmioManager_io_outer_grant_ready),
    .io_outer_grant_valid(mmioManager_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(mmioManager_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(mmioManager_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(mmioManager_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(mmioManager_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(mmioManager_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(mmioManager_io_outer_grant_bits_data)
  );
  Queue_8 Queue_8_1 (
    .clk(Queue_8_1_clk),
    .reset(Queue_8_1_reset),
    .io_enq_ready(Queue_8_1_io_enq_ready),
    .io_enq_valid(Queue_8_1_io_enq_valid),
    .io_enq_bits_addr_block(Queue_8_1_io_enq_bits_addr_block),
    .io_enq_bits_client_xact_id(Queue_8_1_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(Queue_8_1_io_enq_bits_addr_beat),
    .io_enq_bits_is_builtin_type(Queue_8_1_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(Queue_8_1_io_enq_bits_a_type),
    .io_enq_bits_union(Queue_8_1_io_enq_bits_union),
    .io_enq_bits_data(Queue_8_1_io_enq_bits_data),
    .io_deq_ready(Queue_8_1_io_deq_ready),
    .io_deq_valid(Queue_8_1_io_deq_valid),
    .io_deq_bits_addr_block(Queue_8_1_io_deq_bits_addr_block),
    .io_deq_bits_client_xact_id(Queue_8_1_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(Queue_8_1_io_deq_bits_addr_beat),
    .io_deq_bits_is_builtin_type(Queue_8_1_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(Queue_8_1_io_deq_bits_a_type),
    .io_deq_bits_union(Queue_8_1_io_deq_bits_union),
    .io_deq_bits_data(Queue_8_1_io_deq_bits_data),
    .io_count(Queue_8_1_io_count)
  );
  Queue_9 Queue_9_1 (
    .clk(Queue_9_1_clk),
    .reset(Queue_9_1_reset),
    .io_enq_ready(Queue_9_1_io_enq_ready),
    .io_enq_valid(Queue_9_1_io_enq_valid),
    .io_enq_bits_addr_beat(Queue_9_1_io_enq_bits_addr_beat),
    .io_enq_bits_client_xact_id(Queue_9_1_io_enq_bits_client_xact_id),
    .io_enq_bits_manager_xact_id(Queue_9_1_io_enq_bits_manager_xact_id),
    .io_enq_bits_is_builtin_type(Queue_9_1_io_enq_bits_is_builtin_type),
    .io_enq_bits_g_type(Queue_9_1_io_enq_bits_g_type),
    .io_enq_bits_data(Queue_9_1_io_enq_bits_data),
    .io_deq_ready(Queue_9_1_io_deq_ready),
    .io_deq_valid(Queue_9_1_io_deq_valid),
    .io_deq_bits_addr_beat(Queue_9_1_io_deq_bits_addr_beat),
    .io_deq_bits_client_xact_id(Queue_9_1_io_deq_bits_client_xact_id),
    .io_deq_bits_manager_xact_id(Queue_9_1_io_deq_bits_manager_xact_id),
    .io_deq_bits_is_builtin_type(Queue_9_1_io_deq_bits_is_builtin_type),
    .io_deq_bits_g_type(Queue_9_1_io_deq_bits_g_type),
    .io_deq_bits_data(Queue_9_1_io_deq_bits_data),
    .io_count(Queue_9_1_io_count)
  );
  TileLinkMemoryInterconnect mem_ic (
    .clk(mem_ic_clk),
    .reset(mem_ic_reset),
    .io_in_0_acquire_ready(mem_ic_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(mem_ic_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(mem_ic_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(mem_ic_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(mem_ic_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(mem_ic_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(mem_ic_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(mem_ic_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(mem_ic_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(mem_ic_io_in_0_grant_ready),
    .io_in_0_grant_valid(mem_ic_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(mem_ic_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(mem_ic_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(mem_ic_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(mem_ic_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(mem_ic_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(mem_ic_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(mem_ic_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(mem_ic_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(mem_ic_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(mem_ic_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(mem_ic_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(mem_ic_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(mem_ic_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(mem_ic_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(mem_ic_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(mem_ic_io_out_0_grant_ready),
    .io_out_0_grant_valid(mem_ic_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(mem_ic_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(mem_ic_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(mem_ic_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(mem_ic_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(mem_ic_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(mem_ic_io_out_0_grant_bits_data)
  );
  ClientTileLinkIOUnwrapper ClientTileLinkIOUnwrapper_1 (
    .clk(ClientTileLinkIOUnwrapper_1_clk),
    .reset(ClientTileLinkIOUnwrapper_1_reset),
    .io_in_acquire_ready(ClientTileLinkIOUnwrapper_1_io_in_acquire_ready),
    .io_in_acquire_valid(ClientTileLinkIOUnwrapper_1_io_in_acquire_valid),
    .io_in_acquire_bits_addr_block(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_block),
    .io_in_acquire_bits_client_xact_id(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_client_xact_id),
    .io_in_acquire_bits_addr_beat(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_beat),
    .io_in_acquire_bits_is_builtin_type(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_is_builtin_type),
    .io_in_acquire_bits_a_type(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_a_type),
    .io_in_acquire_bits_union(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_union),
    .io_in_acquire_bits_data(ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_data),
    .io_in_probe_ready(ClientTileLinkIOUnwrapper_1_io_in_probe_ready),
    .io_in_probe_valid(ClientTileLinkIOUnwrapper_1_io_in_probe_valid),
    .io_in_probe_bits_addr_block(ClientTileLinkIOUnwrapper_1_io_in_probe_bits_addr_block),
    .io_in_probe_bits_p_type(ClientTileLinkIOUnwrapper_1_io_in_probe_bits_p_type),
    .io_in_release_ready(ClientTileLinkIOUnwrapper_1_io_in_release_ready),
    .io_in_release_valid(ClientTileLinkIOUnwrapper_1_io_in_release_valid),
    .io_in_release_bits_addr_beat(ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_beat),
    .io_in_release_bits_addr_block(ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_block),
    .io_in_release_bits_client_xact_id(ClientTileLinkIOUnwrapper_1_io_in_release_bits_client_xact_id),
    .io_in_release_bits_voluntary(ClientTileLinkIOUnwrapper_1_io_in_release_bits_voluntary),
    .io_in_release_bits_r_type(ClientTileLinkIOUnwrapper_1_io_in_release_bits_r_type),
    .io_in_release_bits_data(ClientTileLinkIOUnwrapper_1_io_in_release_bits_data),
    .io_in_grant_ready(ClientTileLinkIOUnwrapper_1_io_in_grant_ready),
    .io_in_grant_valid(ClientTileLinkIOUnwrapper_1_io_in_grant_valid),
    .io_in_grant_bits_addr_beat(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_addr_beat),
    .io_in_grant_bits_client_xact_id(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_client_xact_id),
    .io_in_grant_bits_manager_xact_id(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_xact_id),
    .io_in_grant_bits_is_builtin_type(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_is_builtin_type),
    .io_in_grant_bits_g_type(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_g_type),
    .io_in_grant_bits_data(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_data),
    .io_in_grant_bits_manager_id(ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_id),
    .io_in_finish_ready(ClientTileLinkIOUnwrapper_1_io_in_finish_ready),
    .io_in_finish_valid(ClientTileLinkIOUnwrapper_1_io_in_finish_valid),
    .io_in_finish_bits_manager_xact_id(ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_xact_id),
    .io_in_finish_bits_manager_id(ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_id),
    .io_out_acquire_ready(ClientTileLinkIOUnwrapper_1_io_out_acquire_ready),
    .io_out_acquire_valid(ClientTileLinkIOUnwrapper_1_io_out_acquire_valid),
    .io_out_acquire_bits_addr_block(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_block),
    .io_out_acquire_bits_client_xact_id(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_client_xact_id),
    .io_out_acquire_bits_addr_beat(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_beat),
    .io_out_acquire_bits_is_builtin_type(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_is_builtin_type),
    .io_out_acquire_bits_a_type(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_a_type),
    .io_out_acquire_bits_union(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_union),
    .io_out_acquire_bits_data(ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_data),
    .io_out_grant_ready(ClientTileLinkIOUnwrapper_1_io_out_grant_ready),
    .io_out_grant_valid(ClientTileLinkIOUnwrapper_1_io_out_grant_valid),
    .io_out_grant_bits_addr_beat(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_addr_beat),
    .io_out_grant_bits_client_xact_id(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_client_xact_id),
    .io_out_grant_bits_manager_xact_id(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_manager_xact_id),
    .io_out_grant_bits_is_builtin_type(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_is_builtin_type),
    .io_out_grant_bits_g_type(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_g_type),
    .io_out_grant_bits_data(ClientTileLinkIOUnwrapper_1_io_out_grant_bits_data)
  );
  ClientTileLinkEnqueuer ClientTileLinkEnqueuer_1 (
    .clk(ClientTileLinkEnqueuer_1_clk),
    .reset(ClientTileLinkEnqueuer_1_reset),
    .io_inner_acquire_ready(ClientTileLinkEnqueuer_1_io_inner_acquire_ready),
    .io_inner_acquire_valid(ClientTileLinkEnqueuer_1_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(ClientTileLinkEnqueuer_1_io_inner_acquire_bits_data),
    .io_inner_probe_ready(ClientTileLinkEnqueuer_1_io_inner_probe_ready),
    .io_inner_probe_valid(ClientTileLinkEnqueuer_1_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(ClientTileLinkEnqueuer_1_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(ClientTileLinkEnqueuer_1_io_inner_probe_bits_p_type),
    .io_inner_release_ready(ClientTileLinkEnqueuer_1_io_inner_release_ready),
    .io_inner_release_valid(ClientTileLinkEnqueuer_1_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(ClientTileLinkEnqueuer_1_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(ClientTileLinkEnqueuer_1_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(ClientTileLinkEnqueuer_1_io_inner_release_bits_data),
    .io_inner_grant_ready(ClientTileLinkEnqueuer_1_io_inner_grant_ready),
    .io_inner_grant_valid(ClientTileLinkEnqueuer_1_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(ClientTileLinkEnqueuer_1_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(ClientTileLinkEnqueuer_1_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(ClientTileLinkEnqueuer_1_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(ClientTileLinkEnqueuer_1_io_inner_grant_bits_data),
    .io_inner_grant_bits_manager_id(ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_id),
    .io_inner_finish_ready(ClientTileLinkEnqueuer_1_io_inner_finish_ready),
    .io_inner_finish_valid(ClientTileLinkEnqueuer_1_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_xact_id),
    .io_inner_finish_bits_manager_id(ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_id),
    .io_outer_acquire_ready(ClientTileLinkEnqueuer_1_io_outer_acquire_ready),
    .io_outer_acquire_valid(ClientTileLinkEnqueuer_1_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(ClientTileLinkEnqueuer_1_io_outer_acquire_bits_data),
    .io_outer_probe_ready(ClientTileLinkEnqueuer_1_io_outer_probe_ready),
    .io_outer_probe_valid(ClientTileLinkEnqueuer_1_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(ClientTileLinkEnqueuer_1_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(ClientTileLinkEnqueuer_1_io_outer_probe_bits_p_type),
    .io_outer_release_ready(ClientTileLinkEnqueuer_1_io_outer_release_ready),
    .io_outer_release_valid(ClientTileLinkEnqueuer_1_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(ClientTileLinkEnqueuer_1_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(ClientTileLinkEnqueuer_1_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(ClientTileLinkEnqueuer_1_io_outer_release_bits_data),
    .io_outer_grant_ready(ClientTileLinkEnqueuer_1_io_outer_grant_ready),
    .io_outer_grant_valid(ClientTileLinkEnqueuer_1_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(ClientTileLinkEnqueuer_1_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(ClientTileLinkEnqueuer_1_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(ClientTileLinkEnqueuer_1_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(ClientTileLinkEnqueuer_1_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(ClientTileLinkEnqueuer_1_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(ClientTileLinkEnqueuer_1_io_outer_finish_ready),
    .io_outer_finish_valid(ClientTileLinkEnqueuer_1_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_id)
  );
  NastiIOTileLinkIOConverter NastiIOTileLinkIOConverter_1 (
    .clk(NastiIOTileLinkIOConverter_1_clk),
    .reset(NastiIOTileLinkIOConverter_1_reset),
    .io_tl_acquire_ready(NastiIOTileLinkIOConverter_1_io_tl_acquire_ready),
    .io_tl_acquire_valid(NastiIOTileLinkIOConverter_1_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_data),
    .io_tl_grant_ready(NastiIOTileLinkIOConverter_1_io_tl_grant_ready),
    .io_tl_grant_valid(NastiIOTileLinkIOConverter_1_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(NastiIOTileLinkIOConverter_1_io_tl_grant_bits_data),
    .io_nasti_aw_ready(NastiIOTileLinkIOConverter_1_io_nasti_aw_ready),
    .io_nasti_aw_valid(NastiIOTileLinkIOConverter_1_io_nasti_aw_valid),
    .io_nasti_aw_bits_addr(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_addr),
    .io_nasti_aw_bits_len(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_len),
    .io_nasti_aw_bits_size(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_size),
    .io_nasti_aw_bits_burst(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_burst),
    .io_nasti_aw_bits_lock(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_lock),
    .io_nasti_aw_bits_cache(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_cache),
    .io_nasti_aw_bits_prot(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_prot),
    .io_nasti_aw_bits_qos(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_qos),
    .io_nasti_aw_bits_region(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_region),
    .io_nasti_aw_bits_id(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_id),
    .io_nasti_aw_bits_user(NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_user),
    .io_nasti_w_ready(NastiIOTileLinkIOConverter_1_io_nasti_w_ready),
    .io_nasti_w_valid(NastiIOTileLinkIOConverter_1_io_nasti_w_valid),
    .io_nasti_w_bits_data(NastiIOTileLinkIOConverter_1_io_nasti_w_bits_data),
    .io_nasti_w_bits_last(NastiIOTileLinkIOConverter_1_io_nasti_w_bits_last),
    .io_nasti_w_bits_id(NastiIOTileLinkIOConverter_1_io_nasti_w_bits_id),
    .io_nasti_w_bits_strb(NastiIOTileLinkIOConverter_1_io_nasti_w_bits_strb),
    .io_nasti_w_bits_user(NastiIOTileLinkIOConverter_1_io_nasti_w_bits_user),
    .io_nasti_b_ready(NastiIOTileLinkIOConverter_1_io_nasti_b_ready),
    .io_nasti_b_valid(NastiIOTileLinkIOConverter_1_io_nasti_b_valid),
    .io_nasti_b_bits_resp(NastiIOTileLinkIOConverter_1_io_nasti_b_bits_resp),
    .io_nasti_b_bits_id(NastiIOTileLinkIOConverter_1_io_nasti_b_bits_id),
    .io_nasti_b_bits_user(NastiIOTileLinkIOConverter_1_io_nasti_b_bits_user),
    .io_nasti_ar_ready(NastiIOTileLinkIOConverter_1_io_nasti_ar_ready),
    .io_nasti_ar_valid(NastiIOTileLinkIOConverter_1_io_nasti_ar_valid),
    .io_nasti_ar_bits_addr(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_addr),
    .io_nasti_ar_bits_len(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_len),
    .io_nasti_ar_bits_size(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_size),
    .io_nasti_ar_bits_burst(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_burst),
    .io_nasti_ar_bits_lock(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_lock),
    .io_nasti_ar_bits_cache(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_cache),
    .io_nasti_ar_bits_prot(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_prot),
    .io_nasti_ar_bits_qos(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_qos),
    .io_nasti_ar_bits_region(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_region),
    .io_nasti_ar_bits_id(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_id),
    .io_nasti_ar_bits_user(NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_user),
    .io_nasti_r_ready(NastiIOTileLinkIOConverter_1_io_nasti_r_ready),
    .io_nasti_r_valid(NastiIOTileLinkIOConverter_1_io_nasti_r_valid),
    .io_nasti_r_bits_resp(NastiIOTileLinkIOConverter_1_io_nasti_r_bits_resp),
    .io_nasti_r_bits_data(NastiIOTileLinkIOConverter_1_io_nasti_r_bits_data),
    .io_nasti_r_bits_last(NastiIOTileLinkIOConverter_1_io_nasti_r_bits_last),
    .io_nasti_r_bits_id(NastiIOTileLinkIOConverter_1_io_nasti_r_bits_id),
    .io_nasti_r_bits_user(NastiIOTileLinkIOConverter_1_io_nasti_r_bits_user)
  );
  Queue_10 Queue_10_1 (
    .clk(Queue_10_1_clk),
    .reset(Queue_10_1_reset),
    .io_enq_ready(Queue_10_1_io_enq_ready),
    .io_enq_valid(Queue_10_1_io_enq_valid),
    .io_enq_bits_addr(Queue_10_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_10_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_10_1_io_enq_bits_size),
    .io_enq_bits_burst(Queue_10_1_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_10_1_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_10_1_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_10_1_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_10_1_io_enq_bits_qos),
    .io_enq_bits_region(Queue_10_1_io_enq_bits_region),
    .io_enq_bits_id(Queue_10_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_10_1_io_enq_bits_user),
    .io_deq_ready(Queue_10_1_io_deq_ready),
    .io_deq_valid(Queue_10_1_io_deq_valid),
    .io_deq_bits_addr(Queue_10_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_10_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_10_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_10_1_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_10_1_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_10_1_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_10_1_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_10_1_io_deq_bits_qos),
    .io_deq_bits_region(Queue_10_1_io_deq_bits_region),
    .io_deq_bits_id(Queue_10_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_10_1_io_deq_bits_user),
    .io_count(Queue_10_1_io_count)
  );
  Queue_10 Queue_11_1 (
    .clk(Queue_11_1_clk),
    .reset(Queue_11_1_reset),
    .io_enq_ready(Queue_11_1_io_enq_ready),
    .io_enq_valid(Queue_11_1_io_enq_valid),
    .io_enq_bits_addr(Queue_11_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_11_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_11_1_io_enq_bits_size),
    .io_enq_bits_burst(Queue_11_1_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_11_1_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_11_1_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_11_1_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_11_1_io_enq_bits_qos),
    .io_enq_bits_region(Queue_11_1_io_enq_bits_region),
    .io_enq_bits_id(Queue_11_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_11_1_io_enq_bits_user),
    .io_deq_ready(Queue_11_1_io_deq_ready),
    .io_deq_valid(Queue_11_1_io_deq_valid),
    .io_deq_bits_addr(Queue_11_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_11_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_11_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_11_1_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_11_1_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_11_1_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_11_1_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_11_1_io_deq_bits_qos),
    .io_deq_bits_region(Queue_11_1_io_deq_bits_region),
    .io_deq_bits_id(Queue_11_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_11_1_io_deq_bits_user),
    .io_count(Queue_11_1_io_count)
  );
  Queue_12 Queue_12_1 (
    .clk(Queue_12_1_clk),
    .reset(Queue_12_1_reset),
    .io_enq_ready(Queue_12_1_io_enq_ready),
    .io_enq_valid(Queue_12_1_io_enq_valid),
    .io_enq_bits_data(Queue_12_1_io_enq_bits_data),
    .io_enq_bits_last(Queue_12_1_io_enq_bits_last),
    .io_enq_bits_id(Queue_12_1_io_enq_bits_id),
    .io_enq_bits_strb(Queue_12_1_io_enq_bits_strb),
    .io_enq_bits_user(Queue_12_1_io_enq_bits_user),
    .io_deq_ready(Queue_12_1_io_deq_ready),
    .io_deq_valid(Queue_12_1_io_deq_valid),
    .io_deq_bits_data(Queue_12_1_io_deq_bits_data),
    .io_deq_bits_last(Queue_12_1_io_deq_bits_last),
    .io_deq_bits_id(Queue_12_1_io_deq_bits_id),
    .io_deq_bits_strb(Queue_12_1_io_deq_bits_strb),
    .io_deq_bits_user(Queue_12_1_io_deq_bits_user),
    .io_count(Queue_12_1_io_count)
  );
  Queue_13 Queue_13_1 (
    .clk(Queue_13_1_clk),
    .reset(Queue_13_1_reset),
    .io_enq_ready(Queue_13_1_io_enq_ready),
    .io_enq_valid(Queue_13_1_io_enq_valid),
    .io_enq_bits_resp(Queue_13_1_io_enq_bits_resp),
    .io_enq_bits_data(Queue_13_1_io_enq_bits_data),
    .io_enq_bits_last(Queue_13_1_io_enq_bits_last),
    .io_enq_bits_id(Queue_13_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_13_1_io_enq_bits_user),
    .io_deq_ready(Queue_13_1_io_deq_ready),
    .io_deq_valid(Queue_13_1_io_deq_valid),
    .io_deq_bits_resp(Queue_13_1_io_deq_bits_resp),
    .io_deq_bits_data(Queue_13_1_io_deq_bits_data),
    .io_deq_bits_last(Queue_13_1_io_deq_bits_last),
    .io_deq_bits_id(Queue_13_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_13_1_io_deq_bits_user),
    .io_count(Queue_13_1_io_count)
  );
  Queue_14 Queue_14_1 (
    .clk(Queue_14_1_clk),
    .reset(Queue_14_1_reset),
    .io_enq_ready(Queue_14_1_io_enq_ready),
    .io_enq_valid(Queue_14_1_io_enq_valid),
    .io_enq_bits_resp(Queue_14_1_io_enq_bits_resp),
    .io_enq_bits_id(Queue_14_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_14_1_io_enq_bits_user),
    .io_deq_ready(Queue_14_1_io_deq_ready),
    .io_deq_valid(Queue_14_1_io_deq_valid),
    .io_deq_bits_resp(Queue_14_1_io_deq_bits_resp),
    .io_deq_bits_id(Queue_14_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_14_1_io_deq_bits_user),
    .io_count(Queue_14_1_io_count)
  );
  assign io_tiles_cached_0_acquire_ready = l1tol2net_io_clients_cached_0_acquire_ready;
  assign io_tiles_cached_0_probe_valid = l1tol2net_io_clients_cached_0_probe_valid;
  assign io_tiles_cached_0_probe_bits_addr_block = l1tol2net_io_clients_cached_0_probe_bits_addr_block;
  assign io_tiles_cached_0_probe_bits_p_type = l1tol2net_io_clients_cached_0_probe_bits_p_type;
  assign io_tiles_cached_0_release_ready = l1tol2net_io_clients_cached_0_release_ready;
  assign io_tiles_cached_0_grant_valid = l1tol2net_io_clients_cached_0_grant_valid;
  assign io_tiles_cached_0_grant_bits_addr_beat = l1tol2net_io_clients_cached_0_grant_bits_addr_beat;
  assign io_tiles_cached_0_grant_bits_client_xact_id = l1tol2net_io_clients_cached_0_grant_bits_client_xact_id;
  assign io_tiles_cached_0_grant_bits_manager_xact_id = l1tol2net_io_clients_cached_0_grant_bits_manager_xact_id;
  assign io_tiles_cached_0_grant_bits_is_builtin_type = l1tol2net_io_clients_cached_0_grant_bits_is_builtin_type;
  assign io_tiles_cached_0_grant_bits_g_type = l1tol2net_io_clients_cached_0_grant_bits_g_type;
  assign io_tiles_cached_0_grant_bits_data = l1tol2net_io_clients_cached_0_grant_bits_data;
  assign io_tiles_cached_0_grant_bits_manager_id = l1tol2net_io_clients_cached_0_grant_bits_manager_id;
  assign io_tiles_cached_0_finish_ready = l1tol2net_io_clients_cached_0_finish_ready;
  assign io_tiles_uncached_0_acquire_ready = l1tol2net_io_clients_uncached_0_acquire_ready;
  assign io_tiles_uncached_0_grant_valid = l1tol2net_io_clients_uncached_0_grant_valid;
  assign io_tiles_uncached_0_grant_bits_addr_beat = l1tol2net_io_clients_uncached_0_grant_bits_addr_beat;
  assign io_tiles_uncached_0_grant_bits_client_xact_id = l1tol2net_io_clients_uncached_0_grant_bits_client_xact_id;
  assign io_tiles_uncached_0_grant_bits_manager_xact_id = l1tol2net_io_clients_uncached_0_grant_bits_manager_xact_id;
  assign io_tiles_uncached_0_grant_bits_is_builtin_type = l1tol2net_io_clients_uncached_0_grant_bits_is_builtin_type;
  assign io_tiles_uncached_0_grant_bits_g_type = l1tol2net_io_clients_uncached_0_grant_bits_g_type;
  assign io_tiles_uncached_0_grant_bits_data = l1tol2net_io_clients_uncached_0_grant_bits_data;
  assign io_mem_axi_0_aw_valid = Queue_11_1_io_deq_valid;
  assign io_mem_axi_0_aw_bits_addr = Queue_11_1_io_deq_bits_addr;
  assign io_mem_axi_0_aw_bits_len = Queue_11_1_io_deq_bits_len;
  assign io_mem_axi_0_aw_bits_size = Queue_11_1_io_deq_bits_size;
  assign io_mem_axi_0_aw_bits_burst = Queue_11_1_io_deq_bits_burst;
  assign io_mem_axi_0_aw_bits_lock = Queue_11_1_io_deq_bits_lock;
  assign io_mem_axi_0_aw_bits_cache = 4'h3;
  assign io_mem_axi_0_aw_bits_prot = Queue_11_1_io_deq_bits_prot;
  assign io_mem_axi_0_aw_bits_qos = Queue_11_1_io_deq_bits_qos;
  assign io_mem_axi_0_aw_bits_region = Queue_11_1_io_deq_bits_region;
  assign io_mem_axi_0_aw_bits_id = Queue_11_1_io_deq_bits_id;
  assign io_mem_axi_0_aw_bits_user = Queue_11_1_io_deq_bits_user;
  assign io_mem_axi_0_w_valid = Queue_12_1_io_deq_valid;
  assign io_mem_axi_0_w_bits_data = Queue_12_1_io_deq_bits_data;
  assign io_mem_axi_0_w_bits_last = Queue_12_1_io_deq_bits_last;
  assign io_mem_axi_0_w_bits_id = Queue_12_1_io_deq_bits_id;
  assign io_mem_axi_0_w_bits_strb = Queue_12_1_io_deq_bits_strb;
  assign io_mem_axi_0_w_bits_user = Queue_12_1_io_deq_bits_user;
  assign io_mem_axi_0_b_ready = Queue_14_1_io_enq_ready;
  assign io_mem_axi_0_ar_valid = Queue_10_1_io_deq_valid;
  assign io_mem_axi_0_ar_bits_addr = Queue_10_1_io_deq_bits_addr;
  assign io_mem_axi_0_ar_bits_len = Queue_10_1_io_deq_bits_len;
  assign io_mem_axi_0_ar_bits_size = Queue_10_1_io_deq_bits_size;
  assign io_mem_axi_0_ar_bits_burst = Queue_10_1_io_deq_bits_burst;
  assign io_mem_axi_0_ar_bits_lock = Queue_10_1_io_deq_bits_lock;
  assign io_mem_axi_0_ar_bits_cache = 4'h3;
  assign io_mem_axi_0_ar_bits_prot = Queue_10_1_io_deq_bits_prot;
  assign io_mem_axi_0_ar_bits_qos = Queue_10_1_io_deq_bits_qos;
  assign io_mem_axi_0_ar_bits_region = Queue_10_1_io_deq_bits_region;
  assign io_mem_axi_0_ar_bits_id = Queue_10_1_io_deq_bits_id;
  assign io_mem_axi_0_ar_bits_user = Queue_10_1_io_deq_bits_user;
  assign io_mem_axi_0_r_ready = Queue_13_1_io_enq_ready;
  assign io_mmio_acquire_valid = Queue_8_1_io_deq_valid;
  assign io_mmio_acquire_bits_addr_block = Queue_8_1_io_deq_bits_addr_block;
  assign io_mmio_acquire_bits_client_xact_id = Queue_8_1_io_deq_bits_client_xact_id;
  assign io_mmio_acquire_bits_addr_beat = Queue_8_1_io_deq_bits_addr_beat;
  assign io_mmio_acquire_bits_is_builtin_type = Queue_8_1_io_deq_bits_is_builtin_type;
  assign io_mmio_acquire_bits_a_type = Queue_8_1_io_deq_bits_a_type;
  assign io_mmio_acquire_bits_union = Queue_8_1_io_deq_bits_union;
  assign io_mmio_acquire_bits_data = Queue_8_1_io_deq_bits_data;
  assign io_mmio_grant_ready = Queue_9_1_io_enq_ready;
  assign l1tol2net_clk = clk;
  assign l1tol2net_reset = reset;
  assign l1tol2net_io_clients_cached_0_acquire_valid = io_tiles_cached_0_acquire_valid;
  assign l1tol2net_io_clients_cached_0_acquire_bits_addr_block = io_tiles_cached_0_acquire_bits_addr_block;
  assign l1tol2net_io_clients_cached_0_acquire_bits_client_xact_id = io_tiles_cached_0_acquire_bits_client_xact_id;
  assign l1tol2net_io_clients_cached_0_acquire_bits_addr_beat = io_tiles_cached_0_acquire_bits_addr_beat;
  assign l1tol2net_io_clients_cached_0_acquire_bits_is_builtin_type = io_tiles_cached_0_acquire_bits_is_builtin_type;
  assign l1tol2net_io_clients_cached_0_acquire_bits_a_type = io_tiles_cached_0_acquire_bits_a_type;
  assign l1tol2net_io_clients_cached_0_acquire_bits_union = io_tiles_cached_0_acquire_bits_union;
  assign l1tol2net_io_clients_cached_0_acquire_bits_data = io_tiles_cached_0_acquire_bits_data;
  assign l1tol2net_io_clients_cached_0_probe_ready = io_tiles_cached_0_probe_ready;
  assign l1tol2net_io_clients_cached_0_release_valid = io_tiles_cached_0_release_valid;
  assign l1tol2net_io_clients_cached_0_release_bits_addr_beat = io_tiles_cached_0_release_bits_addr_beat;
  assign l1tol2net_io_clients_cached_0_release_bits_addr_block = io_tiles_cached_0_release_bits_addr_block;
  assign l1tol2net_io_clients_cached_0_release_bits_client_xact_id = io_tiles_cached_0_release_bits_client_xact_id;
  assign l1tol2net_io_clients_cached_0_release_bits_voluntary = io_tiles_cached_0_release_bits_voluntary;
  assign l1tol2net_io_clients_cached_0_release_bits_r_type = io_tiles_cached_0_release_bits_r_type;
  assign l1tol2net_io_clients_cached_0_release_bits_data = io_tiles_cached_0_release_bits_data;
  assign l1tol2net_io_clients_cached_0_grant_ready = io_tiles_cached_0_grant_ready;
  assign l1tol2net_io_clients_cached_0_finish_valid = io_tiles_cached_0_finish_valid;
  assign l1tol2net_io_clients_cached_0_finish_bits_manager_xact_id = io_tiles_cached_0_finish_bits_manager_xact_id;
  assign l1tol2net_io_clients_cached_0_finish_bits_manager_id = io_tiles_cached_0_finish_bits_manager_id;
  assign l1tol2net_io_clients_uncached_0_acquire_valid = io_tiles_uncached_0_acquire_valid;
  assign l1tol2net_io_clients_uncached_0_acquire_bits_addr_block = io_tiles_uncached_0_acquire_bits_addr_block;
  assign l1tol2net_io_clients_uncached_0_acquire_bits_client_xact_id = io_tiles_uncached_0_acquire_bits_client_xact_id;
  assign l1tol2net_io_clients_uncached_0_acquire_bits_addr_beat = io_tiles_uncached_0_acquire_bits_addr_beat;
  assign l1tol2net_io_clients_uncached_0_acquire_bits_is_builtin_type = io_tiles_uncached_0_acquire_bits_is_builtin_type;
  assign l1tol2net_io_clients_uncached_0_acquire_bits_a_type = io_tiles_uncached_0_acquire_bits_a_type;
  assign l1tol2net_io_clients_uncached_0_acquire_bits_union = io_tiles_uncached_0_acquire_bits_union;
  assign l1tol2net_io_clients_uncached_0_acquire_bits_data = io_tiles_uncached_0_acquire_bits_data;
  assign l1tol2net_io_clients_uncached_0_grant_ready = io_tiles_uncached_0_grant_ready;
  assign l1tol2net_io_managers_0_acquire_ready = ManagerToClientStatelessBridge_1_io_inner_acquire_ready;
  assign l1tol2net_io_managers_0_grant_valid = ManagerToClientStatelessBridge_1_io_inner_grant_valid;
  assign l1tol2net_io_managers_0_grant_bits_addr_beat = ManagerToClientStatelessBridge_1_io_inner_grant_bits_addr_beat;
  assign l1tol2net_io_managers_0_grant_bits_client_xact_id = ManagerToClientStatelessBridge_1_io_inner_grant_bits_client_xact_id;
  assign l1tol2net_io_managers_0_grant_bits_manager_xact_id = ManagerToClientStatelessBridge_1_io_inner_grant_bits_manager_xact_id;
  assign l1tol2net_io_managers_0_grant_bits_is_builtin_type = ManagerToClientStatelessBridge_1_io_inner_grant_bits_is_builtin_type;
  assign l1tol2net_io_managers_0_grant_bits_g_type = ManagerToClientStatelessBridge_1_io_inner_grant_bits_g_type;
  assign l1tol2net_io_managers_0_grant_bits_data = ManagerToClientStatelessBridge_1_io_inner_grant_bits_data;
  assign l1tol2net_io_managers_0_grant_bits_client_id = ManagerToClientStatelessBridge_1_io_inner_grant_bits_client_id;
  assign l1tol2net_io_managers_0_finish_ready = ManagerToClientStatelessBridge_1_io_inner_finish_ready;
  assign l1tol2net_io_managers_0_probe_valid = ManagerToClientStatelessBridge_1_io_inner_probe_valid;
  assign l1tol2net_io_managers_0_probe_bits_addr_block = ManagerToClientStatelessBridge_1_io_inner_probe_bits_addr_block;
  assign l1tol2net_io_managers_0_probe_bits_p_type = ManagerToClientStatelessBridge_1_io_inner_probe_bits_p_type;
  assign l1tol2net_io_managers_0_probe_bits_client_id = ManagerToClientStatelessBridge_1_io_inner_probe_bits_client_id;
  assign l1tol2net_io_managers_0_release_ready = ManagerToClientStatelessBridge_1_io_inner_release_ready;
  assign l1tol2net_io_managers_1_acquire_ready = mmioManager_io_inner_acquire_ready;
  assign l1tol2net_io_managers_1_grant_valid = mmioManager_io_inner_grant_valid;
  assign l1tol2net_io_managers_1_grant_bits_addr_beat = mmioManager_io_inner_grant_bits_addr_beat;
  assign l1tol2net_io_managers_1_grant_bits_client_xact_id = mmioManager_io_inner_grant_bits_client_xact_id;
  assign l1tol2net_io_managers_1_grant_bits_manager_xact_id = mmioManager_io_inner_grant_bits_manager_xact_id;
  assign l1tol2net_io_managers_1_grant_bits_is_builtin_type = mmioManager_io_inner_grant_bits_is_builtin_type;
  assign l1tol2net_io_managers_1_grant_bits_g_type = mmioManager_io_inner_grant_bits_g_type;
  assign l1tol2net_io_managers_1_grant_bits_data = mmioManager_io_inner_grant_bits_data;
  assign l1tol2net_io_managers_1_grant_bits_client_id = mmioManager_io_inner_grant_bits_client_id;
  assign l1tol2net_io_managers_1_finish_ready = mmioManager_io_inner_finish_ready;
  assign l1tol2net_io_managers_1_probe_valid = mmioManager_io_inner_probe_valid;
  assign l1tol2net_io_managers_1_probe_bits_addr_block = mmioManager_io_inner_probe_bits_addr_block;
  assign l1tol2net_io_managers_1_probe_bits_p_type = mmioManager_io_inner_probe_bits_p_type;
  assign l1tol2net_io_managers_1_probe_bits_client_id = mmioManager_io_inner_probe_bits_client_id;
  assign l1tol2net_io_managers_1_release_ready = mmioManager_io_inner_release_ready;
  assign ManagerToClientStatelessBridge_1_clk = clk;
  assign ManagerToClientStatelessBridge_1_reset = reset;
  assign ManagerToClientStatelessBridge_1_io_inner_acquire_valid = l1tol2net_io_managers_0_acquire_valid;
  assign ManagerToClientStatelessBridge_1_io_inner_acquire_bits_addr_block = l1tol2net_io_managers_0_acquire_bits_addr_block;
  assign ManagerToClientStatelessBridge_1_io_inner_acquire_bits_client_xact_id = l1tol2net_io_managers_0_acquire_bits_client_xact_id;
  assign ManagerToClientStatelessBridge_1_io_inner_acquire_bits_addr_beat = l1tol2net_io_managers_0_acquire_bits_addr_beat;
  assign ManagerToClientStatelessBridge_1_io_inner_acquire_bits_is_builtin_type = l1tol2net_io_managers_0_acquire_bits_is_builtin_type;
  assign ManagerToClientStatelessBridge_1_io_inner_acquire_bits_a_type = l1tol2net_io_managers_0_acquire_bits_a_type;
  assign ManagerToClientStatelessBridge_1_io_inner_acquire_bits_union = l1tol2net_io_managers_0_acquire_bits_union;
  assign ManagerToClientStatelessBridge_1_io_inner_acquire_bits_data = l1tol2net_io_managers_0_acquire_bits_data;
  assign ManagerToClientStatelessBridge_1_io_inner_acquire_bits_client_id = l1tol2net_io_managers_0_acquire_bits_client_id;
  assign ManagerToClientStatelessBridge_1_io_inner_grant_ready = l1tol2net_io_managers_0_grant_ready;
  assign ManagerToClientStatelessBridge_1_io_inner_finish_valid = l1tol2net_io_managers_0_finish_valid;
  assign ManagerToClientStatelessBridge_1_io_inner_finish_bits_manager_xact_id = l1tol2net_io_managers_0_finish_bits_manager_xact_id;
  assign ManagerToClientStatelessBridge_1_io_inner_probe_ready = l1tol2net_io_managers_0_probe_ready;
  assign ManagerToClientStatelessBridge_1_io_inner_release_valid = l1tol2net_io_managers_0_release_valid;
  assign ManagerToClientStatelessBridge_1_io_inner_release_bits_addr_beat = l1tol2net_io_managers_0_release_bits_addr_beat;
  assign ManagerToClientStatelessBridge_1_io_inner_release_bits_addr_block = l1tol2net_io_managers_0_release_bits_addr_block;
  assign ManagerToClientStatelessBridge_1_io_inner_release_bits_client_xact_id = l1tol2net_io_managers_0_release_bits_client_xact_id;
  assign ManagerToClientStatelessBridge_1_io_inner_release_bits_voluntary = l1tol2net_io_managers_0_release_bits_voluntary;
  assign ManagerToClientStatelessBridge_1_io_inner_release_bits_r_type = l1tol2net_io_managers_0_release_bits_r_type;
  assign ManagerToClientStatelessBridge_1_io_inner_release_bits_data = l1tol2net_io_managers_0_release_bits_data;
  assign ManagerToClientStatelessBridge_1_io_inner_release_bits_client_id = l1tol2net_io_managers_0_release_bits_client_id;
  assign ManagerToClientStatelessBridge_1_io_incoherent_0 = io_incoherent_0;
  assign ManagerToClientStatelessBridge_1_io_outer_acquire_ready = ClientTileLinkEnqueuer_1_io_inner_acquire_ready;
  assign ManagerToClientStatelessBridge_1_io_outer_probe_valid = ClientTileLinkEnqueuer_1_io_inner_probe_valid;
  assign ManagerToClientStatelessBridge_1_io_outer_probe_bits_addr_block = ClientTileLinkEnqueuer_1_io_inner_probe_bits_addr_block;
  assign ManagerToClientStatelessBridge_1_io_outer_probe_bits_p_type = ClientTileLinkEnqueuer_1_io_inner_probe_bits_p_type;
  assign ManagerToClientStatelessBridge_1_io_outer_release_ready = ClientTileLinkEnqueuer_1_io_inner_release_ready;
  assign ManagerToClientStatelessBridge_1_io_outer_grant_valid = ClientTileLinkEnqueuer_1_io_inner_grant_valid;
  assign ManagerToClientStatelessBridge_1_io_outer_grant_bits_addr_beat = ClientTileLinkEnqueuer_1_io_inner_grant_bits_addr_beat;
  assign ManagerToClientStatelessBridge_1_io_outer_grant_bits_client_xact_id = ClientTileLinkEnqueuer_1_io_inner_grant_bits_client_xact_id;
  assign ManagerToClientStatelessBridge_1_io_outer_grant_bits_manager_xact_id = ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_xact_id;
  assign ManagerToClientStatelessBridge_1_io_outer_grant_bits_is_builtin_type = ClientTileLinkEnqueuer_1_io_inner_grant_bits_is_builtin_type;
  assign ManagerToClientStatelessBridge_1_io_outer_grant_bits_g_type = ClientTileLinkEnqueuer_1_io_inner_grant_bits_g_type;
  assign ManagerToClientStatelessBridge_1_io_outer_grant_bits_data = ClientTileLinkEnqueuer_1_io_inner_grant_bits_data;
  assign ManagerToClientStatelessBridge_1_io_outer_grant_bits_manager_id = ClientTileLinkEnqueuer_1_io_inner_grant_bits_manager_id;
  assign ManagerToClientStatelessBridge_1_io_outer_finish_ready = ClientTileLinkEnqueuer_1_io_inner_finish_ready;
  assign mmioManager_clk = clk;
  assign mmioManager_reset = reset;
  assign mmioManager_io_inner_acquire_valid = l1tol2net_io_managers_1_acquire_valid;
  assign mmioManager_io_inner_acquire_bits_addr_block = l1tol2net_io_managers_1_acquire_bits_addr_block;
  assign mmioManager_io_inner_acquire_bits_client_xact_id = l1tol2net_io_managers_1_acquire_bits_client_xact_id;
  assign mmioManager_io_inner_acquire_bits_addr_beat = l1tol2net_io_managers_1_acquire_bits_addr_beat;
  assign mmioManager_io_inner_acquire_bits_is_builtin_type = l1tol2net_io_managers_1_acquire_bits_is_builtin_type;
  assign mmioManager_io_inner_acquire_bits_a_type = l1tol2net_io_managers_1_acquire_bits_a_type;
  assign mmioManager_io_inner_acquire_bits_union = l1tol2net_io_managers_1_acquire_bits_union;
  assign mmioManager_io_inner_acquire_bits_data = l1tol2net_io_managers_1_acquire_bits_data;
  assign mmioManager_io_inner_acquire_bits_client_id = l1tol2net_io_managers_1_acquire_bits_client_id;
  assign mmioManager_io_inner_grant_ready = l1tol2net_io_managers_1_grant_ready;
  assign mmioManager_io_inner_finish_valid = l1tol2net_io_managers_1_finish_valid;
  assign mmioManager_io_inner_finish_bits_manager_xact_id = l1tol2net_io_managers_1_finish_bits_manager_xact_id;
  assign mmioManager_io_inner_probe_ready = l1tol2net_io_managers_1_probe_ready;
  assign mmioManager_io_inner_release_valid = l1tol2net_io_managers_1_release_valid;
  assign mmioManager_io_inner_release_bits_addr_beat = l1tol2net_io_managers_1_release_bits_addr_beat;
  assign mmioManager_io_inner_release_bits_addr_block = l1tol2net_io_managers_1_release_bits_addr_block;
  assign mmioManager_io_inner_release_bits_client_xact_id = l1tol2net_io_managers_1_release_bits_client_xact_id;
  assign mmioManager_io_inner_release_bits_voluntary = l1tol2net_io_managers_1_release_bits_voluntary;
  assign mmioManager_io_inner_release_bits_r_type = l1tol2net_io_managers_1_release_bits_r_type;
  assign mmioManager_io_inner_release_bits_data = l1tol2net_io_managers_1_release_bits_data;
  assign mmioManager_io_inner_release_bits_client_id = l1tol2net_io_managers_1_release_bits_client_id;
  assign mmioManager_io_incoherent_0 = GEN_0;
  assign mmioManager_io_outer_acquire_ready = Queue_8_1_io_enq_ready;
  assign mmioManager_io_outer_grant_valid = Queue_9_1_io_deq_valid;
  assign mmioManager_io_outer_grant_bits_addr_beat = Queue_9_1_io_deq_bits_addr_beat;
  assign mmioManager_io_outer_grant_bits_client_xact_id = Queue_9_1_io_deq_bits_client_xact_id;
  assign mmioManager_io_outer_grant_bits_manager_xact_id = Queue_9_1_io_deq_bits_manager_xact_id;
  assign mmioManager_io_outer_grant_bits_is_builtin_type = Queue_9_1_io_deq_bits_is_builtin_type;
  assign mmioManager_io_outer_grant_bits_g_type = Queue_9_1_io_deq_bits_g_type;
  assign mmioManager_io_outer_grant_bits_data = Queue_9_1_io_deq_bits_data;
  assign Queue_8_1_clk = clk;
  assign Queue_8_1_reset = reset;
  assign Queue_8_1_io_enq_valid = mmioManager_io_outer_acquire_valid;
  assign Queue_8_1_io_enq_bits_addr_block = mmioManager_io_outer_acquire_bits_addr_block;
  assign Queue_8_1_io_enq_bits_client_xact_id = mmioManager_io_outer_acquire_bits_client_xact_id;
  assign Queue_8_1_io_enq_bits_addr_beat = mmioManager_io_outer_acquire_bits_addr_beat;
  assign Queue_8_1_io_enq_bits_is_builtin_type = mmioManager_io_outer_acquire_bits_is_builtin_type;
  assign Queue_8_1_io_enq_bits_a_type = mmioManager_io_outer_acquire_bits_a_type;
  assign Queue_8_1_io_enq_bits_union = mmioManager_io_outer_acquire_bits_union;
  assign Queue_8_1_io_enq_bits_data = mmioManager_io_outer_acquire_bits_data;
  assign Queue_8_1_io_deq_ready = io_mmio_acquire_ready;
  assign Queue_9_1_clk = clk;
  assign Queue_9_1_reset = reset;
  assign Queue_9_1_io_enq_valid = io_mmio_grant_valid;
  assign Queue_9_1_io_enq_bits_addr_beat = io_mmio_grant_bits_addr_beat;
  assign Queue_9_1_io_enq_bits_client_xact_id = io_mmio_grant_bits_client_xact_id;
  assign Queue_9_1_io_enq_bits_manager_xact_id = io_mmio_grant_bits_manager_xact_id;
  assign Queue_9_1_io_enq_bits_is_builtin_type = io_mmio_grant_bits_is_builtin_type;
  assign Queue_9_1_io_enq_bits_g_type = io_mmio_grant_bits_g_type;
  assign Queue_9_1_io_enq_bits_data = io_mmio_grant_bits_data;
  assign Queue_9_1_io_deq_ready = mmioManager_io_outer_grant_ready;
  assign mem_ic_clk = clk;
  assign mem_ic_reset = reset;
  assign mem_ic_io_in_0_acquire_valid = ClientTileLinkIOUnwrapper_1_io_out_acquire_valid;
  assign mem_ic_io_in_0_acquire_bits_addr_block = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_block;
  assign mem_ic_io_in_0_acquire_bits_client_xact_id = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_client_xact_id;
  assign mem_ic_io_in_0_acquire_bits_addr_beat = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_addr_beat;
  assign mem_ic_io_in_0_acquire_bits_is_builtin_type = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_is_builtin_type;
  assign mem_ic_io_in_0_acquire_bits_a_type = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_a_type;
  assign mem_ic_io_in_0_acquire_bits_union = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_union;
  assign mem_ic_io_in_0_acquire_bits_data = ClientTileLinkIOUnwrapper_1_io_out_acquire_bits_data;
  assign mem_ic_io_in_0_grant_ready = ClientTileLinkIOUnwrapper_1_io_out_grant_ready;
  assign mem_ic_io_out_0_acquire_ready = NastiIOTileLinkIOConverter_1_io_tl_acquire_ready;
  assign mem_ic_io_out_0_grant_valid = NastiIOTileLinkIOConverter_1_io_tl_grant_valid;
  assign mem_ic_io_out_0_grant_bits_addr_beat = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_addr_beat;
  assign mem_ic_io_out_0_grant_bits_client_xact_id = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_client_xact_id;
  assign mem_ic_io_out_0_grant_bits_manager_xact_id = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_manager_xact_id;
  assign mem_ic_io_out_0_grant_bits_is_builtin_type = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_is_builtin_type;
  assign mem_ic_io_out_0_grant_bits_g_type = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_g_type;
  assign mem_ic_io_out_0_grant_bits_data = NastiIOTileLinkIOConverter_1_io_tl_grant_bits_data;
  assign ClientTileLinkIOUnwrapper_1_clk = clk;
  assign ClientTileLinkIOUnwrapper_1_reset = reset;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_valid = ClientTileLinkEnqueuer_1_io_outer_acquire_valid;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_block = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_block;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_client_xact_id = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_client_xact_id;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_addr_beat = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_addr_beat;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_is_builtin_type = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_is_builtin_type;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_a_type = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_a_type;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_union = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_union;
  assign ClientTileLinkIOUnwrapper_1_io_in_acquire_bits_data = ClientTileLinkEnqueuer_1_io_outer_acquire_bits_data;
  assign ClientTileLinkIOUnwrapper_1_io_in_probe_ready = ClientTileLinkEnqueuer_1_io_outer_probe_ready;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_valid = ClientTileLinkEnqueuer_1_io_outer_release_valid;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_beat = ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_beat;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_addr_block = ClientTileLinkEnqueuer_1_io_outer_release_bits_addr_block;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_client_xact_id = ClientTileLinkEnqueuer_1_io_outer_release_bits_client_xact_id;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_voluntary = ClientTileLinkEnqueuer_1_io_outer_release_bits_voluntary;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_r_type = ClientTileLinkEnqueuer_1_io_outer_release_bits_r_type;
  assign ClientTileLinkIOUnwrapper_1_io_in_release_bits_data = ClientTileLinkEnqueuer_1_io_outer_release_bits_data;
  assign ClientTileLinkIOUnwrapper_1_io_in_grant_ready = ClientTileLinkEnqueuer_1_io_outer_grant_ready;
  assign ClientTileLinkIOUnwrapper_1_io_in_finish_valid = ClientTileLinkEnqueuer_1_io_outer_finish_valid;
  assign ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_xact_id = ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_xact_id;
  assign ClientTileLinkIOUnwrapper_1_io_in_finish_bits_manager_id = ClientTileLinkEnqueuer_1_io_outer_finish_bits_manager_id;
  assign ClientTileLinkIOUnwrapper_1_io_out_acquire_ready = mem_ic_io_in_0_acquire_ready;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_valid = mem_ic_io_in_0_grant_valid;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_addr_beat = mem_ic_io_in_0_grant_bits_addr_beat;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_client_xact_id = mem_ic_io_in_0_grant_bits_client_xact_id;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_manager_xact_id = mem_ic_io_in_0_grant_bits_manager_xact_id;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_is_builtin_type = mem_ic_io_in_0_grant_bits_is_builtin_type;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_g_type = mem_ic_io_in_0_grant_bits_g_type;
  assign ClientTileLinkIOUnwrapper_1_io_out_grant_bits_data = mem_ic_io_in_0_grant_bits_data;
  assign ClientTileLinkEnqueuer_1_clk = clk;
  assign ClientTileLinkEnqueuer_1_reset = reset;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_valid = ManagerToClientStatelessBridge_1_io_outer_acquire_valid;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_block = ManagerToClientStatelessBridge_1_io_outer_acquire_bits_addr_block;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_client_xact_id = ManagerToClientStatelessBridge_1_io_outer_acquire_bits_client_xact_id;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_addr_beat = ManagerToClientStatelessBridge_1_io_outer_acquire_bits_addr_beat;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_is_builtin_type = ManagerToClientStatelessBridge_1_io_outer_acquire_bits_is_builtin_type;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_a_type = ManagerToClientStatelessBridge_1_io_outer_acquire_bits_a_type;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_union = ManagerToClientStatelessBridge_1_io_outer_acquire_bits_union;
  assign ClientTileLinkEnqueuer_1_io_inner_acquire_bits_data = ManagerToClientStatelessBridge_1_io_outer_acquire_bits_data;
  assign ClientTileLinkEnqueuer_1_io_inner_probe_ready = ManagerToClientStatelessBridge_1_io_outer_probe_ready;
  assign ClientTileLinkEnqueuer_1_io_inner_release_valid = ManagerToClientStatelessBridge_1_io_outer_release_valid;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_beat = ManagerToClientStatelessBridge_1_io_outer_release_bits_addr_beat;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_addr_block = ManagerToClientStatelessBridge_1_io_outer_release_bits_addr_block;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_client_xact_id = ManagerToClientStatelessBridge_1_io_outer_release_bits_client_xact_id;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_voluntary = ManagerToClientStatelessBridge_1_io_outer_release_bits_voluntary;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_r_type = ManagerToClientStatelessBridge_1_io_outer_release_bits_r_type;
  assign ClientTileLinkEnqueuer_1_io_inner_release_bits_data = ManagerToClientStatelessBridge_1_io_outer_release_bits_data;
  assign ClientTileLinkEnqueuer_1_io_inner_grant_ready = ManagerToClientStatelessBridge_1_io_outer_grant_ready;
  assign ClientTileLinkEnqueuer_1_io_inner_finish_valid = ManagerToClientStatelessBridge_1_io_outer_finish_valid;
  assign ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_xact_id = ManagerToClientStatelessBridge_1_io_outer_finish_bits_manager_xact_id;
  assign ClientTileLinkEnqueuer_1_io_inner_finish_bits_manager_id = ManagerToClientStatelessBridge_1_io_outer_finish_bits_manager_id;
  assign ClientTileLinkEnqueuer_1_io_outer_acquire_ready = ClientTileLinkIOUnwrapper_1_io_in_acquire_ready;
  assign ClientTileLinkEnqueuer_1_io_outer_probe_valid = ClientTileLinkIOUnwrapper_1_io_in_probe_valid;
  assign ClientTileLinkEnqueuer_1_io_outer_probe_bits_addr_block = ClientTileLinkIOUnwrapper_1_io_in_probe_bits_addr_block;
  assign ClientTileLinkEnqueuer_1_io_outer_probe_bits_p_type = ClientTileLinkIOUnwrapper_1_io_in_probe_bits_p_type;
  assign ClientTileLinkEnqueuer_1_io_outer_release_ready = ClientTileLinkIOUnwrapper_1_io_in_release_ready;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_valid = ClientTileLinkIOUnwrapper_1_io_in_grant_valid;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_addr_beat = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_addr_beat;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_client_xact_id = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_client_xact_id;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_xact_id = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_xact_id;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_is_builtin_type = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_is_builtin_type;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_g_type = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_g_type;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_data = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_data;
  assign ClientTileLinkEnqueuer_1_io_outer_grant_bits_manager_id = ClientTileLinkIOUnwrapper_1_io_in_grant_bits_manager_id;
  assign ClientTileLinkEnqueuer_1_io_outer_finish_ready = ClientTileLinkIOUnwrapper_1_io_in_finish_ready;
  assign NastiIOTileLinkIOConverter_1_clk = clk;
  assign NastiIOTileLinkIOConverter_1_reset = reset;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_valid = mem_ic_io_out_0_acquire_valid;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_block = mem_ic_io_out_0_acquire_bits_addr_block;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_client_xact_id = mem_ic_io_out_0_acquire_bits_client_xact_id;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_addr_beat = mem_ic_io_out_0_acquire_bits_addr_beat;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_is_builtin_type = mem_ic_io_out_0_acquire_bits_is_builtin_type;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_a_type = mem_ic_io_out_0_acquire_bits_a_type;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_union = mem_ic_io_out_0_acquire_bits_union;
  assign NastiIOTileLinkIOConverter_1_io_tl_acquire_bits_data = mem_ic_io_out_0_acquire_bits_data;
  assign NastiIOTileLinkIOConverter_1_io_tl_grant_ready = mem_ic_io_out_0_grant_ready;
  assign NastiIOTileLinkIOConverter_1_io_nasti_aw_ready = Queue_11_1_io_enq_ready;
  assign NastiIOTileLinkIOConverter_1_io_nasti_w_ready = Queue_12_1_io_enq_ready;
  assign NastiIOTileLinkIOConverter_1_io_nasti_b_valid = Queue_14_1_io_deq_valid;
  assign NastiIOTileLinkIOConverter_1_io_nasti_b_bits_resp = Queue_14_1_io_deq_bits_resp;
  assign NastiIOTileLinkIOConverter_1_io_nasti_b_bits_id = Queue_14_1_io_deq_bits_id;
  assign NastiIOTileLinkIOConverter_1_io_nasti_b_bits_user = Queue_14_1_io_deq_bits_user;
  assign NastiIOTileLinkIOConverter_1_io_nasti_ar_ready = Queue_10_1_io_enq_ready;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_valid = Queue_13_1_io_deq_valid;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_bits_resp = Queue_13_1_io_deq_bits_resp;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_bits_data = Queue_13_1_io_deq_bits_data;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_bits_last = Queue_13_1_io_deq_bits_last;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_bits_id = Queue_13_1_io_deq_bits_id;
  assign NastiIOTileLinkIOConverter_1_io_nasti_r_bits_user = Queue_13_1_io_deq_bits_user;
  assign Queue_10_1_clk = clk;
  assign Queue_10_1_reset = reset;
  assign Queue_10_1_io_enq_valid = NastiIOTileLinkIOConverter_1_io_nasti_ar_valid;
  assign Queue_10_1_io_enq_bits_addr = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_addr;
  assign Queue_10_1_io_enq_bits_len = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_len;
  assign Queue_10_1_io_enq_bits_size = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_size;
  assign Queue_10_1_io_enq_bits_burst = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_burst;
  assign Queue_10_1_io_enq_bits_lock = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_lock;
  assign Queue_10_1_io_enq_bits_cache = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_cache;
  assign Queue_10_1_io_enq_bits_prot = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_prot;
  assign Queue_10_1_io_enq_bits_qos = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_qos;
  assign Queue_10_1_io_enq_bits_region = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_region;
  assign Queue_10_1_io_enq_bits_id = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_id;
  assign Queue_10_1_io_enq_bits_user = NastiIOTileLinkIOConverter_1_io_nasti_ar_bits_user;
  assign Queue_10_1_io_deq_ready = io_mem_axi_0_ar_ready;
  assign Queue_11_1_clk = clk;
  assign Queue_11_1_reset = reset;
  assign Queue_11_1_io_enq_valid = NastiIOTileLinkIOConverter_1_io_nasti_aw_valid;
  assign Queue_11_1_io_enq_bits_addr = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_addr;
  assign Queue_11_1_io_enq_bits_len = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_len;
  assign Queue_11_1_io_enq_bits_size = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_size;
  assign Queue_11_1_io_enq_bits_burst = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_burst;
  assign Queue_11_1_io_enq_bits_lock = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_lock;
  assign Queue_11_1_io_enq_bits_cache = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_cache;
  assign Queue_11_1_io_enq_bits_prot = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_prot;
  assign Queue_11_1_io_enq_bits_qos = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_qos;
  assign Queue_11_1_io_enq_bits_region = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_region;
  assign Queue_11_1_io_enq_bits_id = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_id;
  assign Queue_11_1_io_enq_bits_user = NastiIOTileLinkIOConverter_1_io_nasti_aw_bits_user;
  assign Queue_11_1_io_deq_ready = io_mem_axi_0_aw_ready;
  assign Queue_12_1_clk = clk;
  assign Queue_12_1_reset = reset;
  assign Queue_12_1_io_enq_valid = NastiIOTileLinkIOConverter_1_io_nasti_w_valid;
  assign Queue_12_1_io_enq_bits_data = NastiIOTileLinkIOConverter_1_io_nasti_w_bits_data;
  assign Queue_12_1_io_enq_bits_last = NastiIOTileLinkIOConverter_1_io_nasti_w_bits_last;
  assign Queue_12_1_io_enq_bits_id = NastiIOTileLinkIOConverter_1_io_nasti_w_bits_id;
  assign Queue_12_1_io_enq_bits_strb = NastiIOTileLinkIOConverter_1_io_nasti_w_bits_strb;
  assign Queue_12_1_io_enq_bits_user = NastiIOTileLinkIOConverter_1_io_nasti_w_bits_user;
  assign Queue_12_1_io_deq_ready = io_mem_axi_0_w_ready;
  assign Queue_13_1_clk = clk;
  assign Queue_13_1_reset = reset;
  assign Queue_13_1_io_enq_valid = io_mem_axi_0_r_valid;
  assign Queue_13_1_io_enq_bits_resp = io_mem_axi_0_r_bits_resp;
  assign Queue_13_1_io_enq_bits_data = io_mem_axi_0_r_bits_data;
  assign Queue_13_1_io_enq_bits_last = io_mem_axi_0_r_bits_last;
  assign Queue_13_1_io_enq_bits_id = io_mem_axi_0_r_bits_id;
  assign Queue_13_1_io_enq_bits_user = io_mem_axi_0_r_bits_user;
  assign Queue_13_1_io_deq_ready = NastiIOTileLinkIOConverter_1_io_nasti_r_ready;
  assign Queue_14_1_clk = clk;
  assign Queue_14_1_reset = reset;
  assign Queue_14_1_io_enq_valid = io_mem_axi_0_b_valid;
  assign Queue_14_1_io_enq_bits_resp = io_mem_axi_0_b_bits_resp;
  assign Queue_14_1_io_enq_bits_id = io_mem_axi_0_b_bits_id;
  assign Queue_14_1_io_enq_bits_user = io_mem_axi_0_b_bits_user;
  assign Queue_14_1_io_deq_ready = NastiIOTileLinkIOConverter_1_io_nasti_b_ready;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_1 = {1{$random}};
  GEN_0 = GEN_1[0:0];
  `endif
  end
`endif
endmodule
module LockingRRArbiter_6(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [1:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_is_builtin_type,
  input  [3:0] io_in_1_bits_g_type,
  input  [63:0] io_in_1_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_chosen
);
  wire  choice;
  wire  GEN_0;
  wire  GEN_7;
  wire [2:0] GEN_1;
  wire [2:0] GEN_8;
  wire [1:0] GEN_2;
  wire [1:0] GEN_9;
  wire  GEN_3;
  wire  GEN_10;
  wire  GEN_4;
  wire  GEN_11;
  wire [3:0] GEN_5;
  wire [3:0] GEN_12;
  wire [63:0] GEN_6;
  wire [63:0] GEN_13;
  reg [2:0] T_610;
  reg [31:0] GEN_21;
  reg  T_612;
  reg [31:0] GEN_22;
  wire  T_614;
  wire [2:0] T_622_0;
  wire [3:0] GEN_20;
  wire  T_624;
  wire  T_625;
  wire  T_626;
  wire  T_628;
  wire  T_629;
  wire [3:0] T_633;
  wire [2:0] T_634;
  wire  GEN_14;
  wire [2:0] GEN_15;
  wire  GEN_16;
  reg  lastGrant;
  reg [31:0] GEN_23;
  wire  GEN_17;
  wire  T_639;
  wire  T_641;
  wire  T_644;
  wire  T_648;
  wire  T_650;
  wire  T_654;
  wire  T_656;
  wire  T_657;
  wire  T_658;
  wire  T_661;
  wire  T_662;
  wire  GEN_18;
  wire  GEN_19;
  assign io_in_0_ready = T_658;
  assign io_in_1_ready = T_662;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_beat = GEN_1;
  assign io_out_bits_client_xact_id = GEN_2;
  assign io_out_bits_manager_xact_id = GEN_3;
  assign io_out_bits_is_builtin_type = GEN_4;
  assign io_out_bits_g_type = GEN_5;
  assign io_out_bits_data = GEN_6;
  assign io_chosen = GEN_16;
  assign choice = GEN_19;
  assign GEN_0 = GEN_7;
  assign GEN_7 = io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_1 = GEN_8;
  assign GEN_8 = io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_2 = GEN_9;
  assign GEN_9 = io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_3 = GEN_10;
  assign GEN_10 = io_chosen ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign GEN_4 = GEN_11;
  assign GEN_11 = io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_5 = GEN_12;
  assign GEN_12 = io_chosen ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign GEN_6 = GEN_13;
  assign GEN_13 = io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign T_614 = T_610 != 3'h0;
  assign T_622_0 = 3'h5;
  assign GEN_20 = {{1'd0}, T_622_0};
  assign T_624 = io_out_bits_g_type == GEN_20;
  assign T_625 = io_out_bits_g_type == 4'h0;
  assign T_626 = io_out_bits_is_builtin_type ? T_624 : T_625;
  assign T_628 = io_out_ready & io_out_valid;
  assign T_629 = T_628 & T_626;
  assign T_633 = T_610 + 3'h1;
  assign T_634 = T_633[2:0];
  assign GEN_14 = T_629 ? io_chosen : T_612;
  assign GEN_15 = T_629 ? T_634 : T_610;
  assign GEN_16 = T_614 ? T_612 : choice;
  assign GEN_17 = T_628 ? io_chosen : lastGrant;
  assign T_639 = 1'h1 > lastGrant;
  assign T_641 = io_in_1_valid & T_639;
  assign T_644 = T_641 | io_in_0_valid;
  assign T_648 = T_641 == 1'h0;
  assign T_650 = T_644 == 1'h0;
  assign T_654 = T_639 | T_650;
  assign T_656 = T_612 == 1'h0;
  assign T_657 = T_614 ? T_656 : T_648;
  assign T_658 = T_657 & io_out_ready;
  assign T_661 = T_614 ? T_612 : T_654;
  assign T_662 = T_661 & io_out_ready;
  assign GEN_18 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_19 = T_641 ? 1'h1 : GEN_18;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_21 = {1{$random}};
  T_610 = GEN_21[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_22 = {1{$random}};
  T_612 = GEN_22[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_23 = {1{$random}};
  lastGrant = GEN_23[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_610 <= 3'h0;
    end else begin
      if(T_629) begin
        T_610 <= T_634;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_629) begin
        T_612 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_628) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module ClientUncachedTileLinkIORouter(
  input   clk,
  input   reset,
  output  io_in_acquire_ready,
  input   io_in_acquire_valid,
  input  [25:0] io_in_acquire_bits_addr_block,
  input  [1:0] io_in_acquire_bits_client_xact_id,
  input  [2:0] io_in_acquire_bits_addr_beat,
  input   io_in_acquire_bits_is_builtin_type,
  input  [2:0] io_in_acquire_bits_a_type,
  input  [11:0] io_in_acquire_bits_union,
  input  [63:0] io_in_acquire_bits_data,
  input   io_in_grant_ready,
  output  io_in_grant_valid,
  output [2:0] io_in_grant_bits_addr_beat,
  output [1:0] io_in_grant_bits_client_xact_id,
  output  io_in_grant_bits_manager_xact_id,
  output  io_in_grant_bits_is_builtin_type,
  output [3:0] io_in_grant_bits_g_type,
  output [63:0] io_in_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [11:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [11:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data
);
  wire [2:0] T_1449_0;
  wire [2:0] T_1449_1;
  wire  T_1451;
  wire  T_1452;
  wire  T_1453;
  wire  T_1454;
  wire [2:0] T_1455;
  wire [2:0] T_1457;
  wire [28:0] T_1458;
  wire [31:0] T_1459;
  wire  T_1463;
  wire  T_1466;
  wire  T_1468;
  wire  T_1469;
  wire [1:0] acq_route;
  wire  T_1471;
  wire  T_1472;
  wire  GEN_0;
  wire  T_1474;
  wire  T_1475;
  wire  GEN_1;
  wire  gnt_arb_clk;
  wire  gnt_arb_reset;
  wire  gnt_arb_io_in_0_ready;
  wire  gnt_arb_io_in_0_valid;
  wire [2:0] gnt_arb_io_in_0_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_0_bits_client_xact_id;
  wire  gnt_arb_io_in_0_bits_manager_xact_id;
  wire  gnt_arb_io_in_0_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_0_bits_g_type;
  wire [63:0] gnt_arb_io_in_0_bits_data;
  wire  gnt_arb_io_in_1_ready;
  wire  gnt_arb_io_in_1_valid;
  wire [2:0] gnt_arb_io_in_1_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_1_bits_client_xact_id;
  wire  gnt_arb_io_in_1_bits_manager_xact_id;
  wire  gnt_arb_io_in_1_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_1_bits_g_type;
  wire [63:0] gnt_arb_io_in_1_bits_data;
  wire  gnt_arb_io_out_ready;
  wire  gnt_arb_io_out_valid;
  wire [2:0] gnt_arb_io_out_bits_addr_beat;
  wire [1:0] gnt_arb_io_out_bits_client_xact_id;
  wire  gnt_arb_io_out_bits_manager_xact_id;
  wire  gnt_arb_io_out_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_out_bits_g_type;
  wire [63:0] gnt_arb_io_out_bits_data;
  wire  gnt_arb_io_chosen;
  wire  T_1500;
  wire  T_1502;
  wire  T_1503;
  wire  T_1504;
  wire  T_1506;
  LockingRRArbiter_6 gnt_arb (
    .clk(gnt_arb_clk),
    .reset(gnt_arb_reset),
    .io_in_0_ready(gnt_arb_io_in_0_ready),
    .io_in_0_valid(gnt_arb_io_in_0_valid),
    .io_in_0_bits_addr_beat(gnt_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(gnt_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(gnt_arb_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(gnt_arb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(gnt_arb_io_in_0_bits_g_type),
    .io_in_0_bits_data(gnt_arb_io_in_0_bits_data),
    .io_in_1_ready(gnt_arb_io_in_1_ready),
    .io_in_1_valid(gnt_arb_io_in_1_valid),
    .io_in_1_bits_addr_beat(gnt_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_client_xact_id(gnt_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_manager_xact_id(gnt_arb_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_is_builtin_type(gnt_arb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_g_type(gnt_arb_io_in_1_bits_g_type),
    .io_in_1_bits_data(gnt_arb_io_in_1_bits_data),
    .io_out_ready(gnt_arb_io_out_ready),
    .io_out_valid(gnt_arb_io_out_valid),
    .io_out_bits_addr_beat(gnt_arb_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(gnt_arb_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(gnt_arb_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(gnt_arb_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(gnt_arb_io_out_bits_g_type),
    .io_out_bits_data(gnt_arb_io_out_bits_data),
    .io_chosen(gnt_arb_io_chosen)
  );
  assign io_in_acquire_ready = GEN_1;
  assign io_in_grant_valid = gnt_arb_io_out_valid;
  assign io_in_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_in_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_in_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_in_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_in_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_in_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_out_0_acquire_valid = T_1472;
  assign io_out_0_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_0_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_0_grant_ready = gnt_arb_io_in_0_ready;
  assign io_out_1_acquire_valid = T_1475;
  assign io_out_1_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_1_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_1_grant_ready = gnt_arb_io_in_1_ready;
  assign T_1449_0 = 3'h0;
  assign T_1449_1 = 3'h4;
  assign T_1451 = io_in_acquire_bits_a_type == T_1449_0;
  assign T_1452 = io_in_acquire_bits_a_type == T_1449_1;
  assign T_1453 = T_1451 | T_1452;
  assign T_1454 = io_in_acquire_bits_is_builtin_type & T_1453;
  assign T_1455 = io_in_acquire_bits_union[11:9];
  assign T_1457 = T_1454 ? T_1455 : 3'h0;
  assign T_1458 = {io_in_acquire_bits_addr_block,io_in_acquire_bits_addr_beat};
  assign T_1459 = {T_1458,T_1457};
  assign T_1463 = T_1459 < 32'h48000000;
  assign T_1466 = 32'h60000000 <= T_1459;
  assign T_1468 = T_1459 < 32'h80000000;
  assign T_1469 = T_1466 & T_1468;
  assign acq_route = {T_1469,T_1463};
  assign T_1471 = acq_route[0];
  assign T_1472 = io_in_acquire_valid & T_1471;
  assign GEN_0 = T_1471 ? io_out_0_acquire_ready : 1'h0;
  assign T_1474 = acq_route[1];
  assign T_1475 = io_in_acquire_valid & T_1474;
  assign GEN_1 = T_1474 ? io_out_1_acquire_ready : GEN_0;
  assign gnt_arb_clk = clk;
  assign gnt_arb_reset = reset;
  assign gnt_arb_io_in_0_valid = io_out_0_grant_valid;
  assign gnt_arb_io_in_0_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign gnt_arb_io_in_0_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign gnt_arb_io_in_0_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_0_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_0_bits_g_type = io_out_0_grant_bits_g_type;
  assign gnt_arb_io_in_0_bits_data = io_out_0_grant_bits_data;
  assign gnt_arb_io_in_1_valid = io_out_1_grant_valid;
  assign gnt_arb_io_in_1_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign gnt_arb_io_in_1_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign gnt_arb_io_in_1_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_1_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_1_bits_g_type = io_out_1_grant_bits_g_type;
  assign gnt_arb_io_in_1_bits_data = io_out_1_grant_bits_data;
  assign gnt_arb_io_out_ready = io_in_grant_ready;
  assign T_1500 = io_in_acquire_valid == 1'h0;
  assign T_1502 = acq_route != 2'h0;
  assign T_1503 = T_1500 | T_1502;
  assign T_1504 = T_1503 | reset;
  assign T_1506 = T_1504 == 1'h0;
  always @(posedge clk) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1506) begin
          $fwrite(32'h80000002,"Assertion failed: No valid route\n    at Interconnect.scala:219 assert(!io.in.acquire.valid || acq_route.orR, ---No valid route---)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1506) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module ClientUncachedTileLinkIOCrossbar(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [11:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [11:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data
);
  wire  ClientUncachedTileLinkIORouter_1_clk;
  wire  ClientUncachedTileLinkIORouter_1_reset;
  wire  ClientUncachedTileLinkIORouter_1_io_in_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_io_in_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_io_in_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_io_in_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_in_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_io_in_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_io_in_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_io_in_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_io_in_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_io_in_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_io_out_1_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_io_out_1_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_io_out_1_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_io_out_1_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_data;
  ClientUncachedTileLinkIORouter ClientUncachedTileLinkIORouter_1 (
    .clk(ClientUncachedTileLinkIORouter_1_clk),
    .reset(ClientUncachedTileLinkIORouter_1_reset),
    .io_in_acquire_ready(ClientUncachedTileLinkIORouter_1_io_in_acquire_ready),
    .io_in_acquire_valid(ClientUncachedTileLinkIORouter_1_io_in_acquire_valid),
    .io_in_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_block),
    .io_in_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_client_xact_id),
    .io_in_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_beat),
    .io_in_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_is_builtin_type),
    .io_in_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_a_type),
    .io_in_acquire_bits_union(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_union),
    .io_in_acquire_bits_data(ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_data),
    .io_in_grant_ready(ClientUncachedTileLinkIORouter_1_io_in_grant_ready),
    .io_in_grant_valid(ClientUncachedTileLinkIORouter_1_io_in_grant_valid),
    .io_in_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_addr_beat),
    .io_in_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_client_xact_id),
    .io_in_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_manager_xact_id),
    .io_in_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_is_builtin_type),
    .io_in_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_g_type),
    .io_in_grant_bits_data(ClientUncachedTileLinkIORouter_1_io_in_grant_bits_data),
    .io_out_0_acquire_ready(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(ClientUncachedTileLinkIORouter_1_io_out_0_grant_ready),
    .io_out_0_grant_valid(ClientUncachedTileLinkIORouter_1_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(ClientUncachedTileLinkIORouter_1_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(ClientUncachedTileLinkIORouter_1_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(ClientUncachedTileLinkIORouter_1_io_out_1_grant_ready),
    .io_out_1_grant_valid(ClientUncachedTileLinkIORouter_1_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_data)
  );
  assign io_in_0_acquire_ready = ClientUncachedTileLinkIORouter_1_io_in_acquire_ready;
  assign io_in_0_grant_valid = ClientUncachedTileLinkIORouter_1_io_in_grant_valid;
  assign io_in_0_grant_bits_addr_beat = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_g_type;
  assign io_in_0_grant_bits_data = ClientUncachedTileLinkIORouter_1_io_in_grant_bits_data;
  assign io_out_0_acquire_valid = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_union;
  assign io_out_0_acquire_bits_data = ClientUncachedTileLinkIORouter_1_io_out_0_acquire_bits_data;
  assign io_out_0_grant_ready = ClientUncachedTileLinkIORouter_1_io_out_0_grant_ready;
  assign io_out_1_acquire_valid = ClientUncachedTileLinkIORouter_1_io_out_1_acquire_valid;
  assign io_out_1_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_union;
  assign io_out_1_acquire_bits_data = ClientUncachedTileLinkIORouter_1_io_out_1_acquire_bits_data;
  assign io_out_1_grant_ready = ClientUncachedTileLinkIORouter_1_io_out_1_grant_ready;
  assign ClientUncachedTileLinkIORouter_1_clk = clk;
  assign ClientUncachedTileLinkIORouter_1_reset = reset;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_valid = io_in_0_acquire_valid;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_union = io_in_0_acquire_bits_union;
  assign ClientUncachedTileLinkIORouter_1_io_in_acquire_bits_data = io_in_0_acquire_bits_data;
  assign ClientUncachedTileLinkIORouter_1_io_in_grant_ready = io_in_0_grant_ready;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_acquire_ready = io_out_0_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_valid = io_out_0_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_io_out_0_grant_bits_data = io_out_0_grant_bits_data;
  assign ClientUncachedTileLinkIORouter_1_io_out_1_acquire_ready = io_out_1_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_io_out_1_grant_valid = io_out_1_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_g_type = io_out_1_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_io_out_1_grant_bits_data = io_out_1_grant_bits_data;
endmodule
module LockingRRArbiter_7(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [1:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_is_builtin_type,
  input  [3:0] io_in_1_bits_g_type,
  input  [63:0] io_in_1_bits_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_addr_beat,
  input  [1:0] io_in_2_bits_client_xact_id,
  input   io_in_2_bits_manager_xact_id,
  input   io_in_2_bits_is_builtin_type,
  input  [3:0] io_in_2_bits_g_type,
  input  [63:0] io_in_2_bits_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [2:0] io_in_3_bits_addr_beat,
  input  [1:0] io_in_3_bits_client_xact_id,
  input   io_in_3_bits_manager_xact_id,
  input   io_in_3_bits_is_builtin_type,
  input  [3:0] io_in_3_bits_g_type,
  input  [63:0] io_in_3_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire [2:0] GEN_1;
  wire [2:0] GEN_10;
  wire [2:0] GEN_11;
  wire [2:0] GEN_12;
  wire [1:0] GEN_2;
  wire [1:0] GEN_13;
  wire [1:0] GEN_14;
  wire [1:0] GEN_15;
  wire  GEN_3;
  wire  GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire  GEN_4;
  wire  GEN_19;
  wire  GEN_20;
  wire  GEN_21;
  wire [3:0] GEN_5;
  wire [3:0] GEN_22;
  wire [3:0] GEN_23;
  wire [3:0] GEN_24;
  wire [63:0] GEN_6;
  wire [63:0] GEN_25;
  wire [63:0] GEN_26;
  wire [63:0] GEN_27;
  reg [2:0] T_794;
  reg [31:0] GEN_39;
  reg [1:0] T_796;
  reg [31:0] GEN_40;
  wire  T_798;
  wire [2:0] T_806_0;
  wire [3:0] GEN_38;
  wire  T_808;
  wire  T_809;
  wire  T_810;
  wire  T_812;
  wire  T_813;
  wire [3:0] T_817;
  wire [2:0] T_818;
  wire [1:0] GEN_28;
  wire [2:0] GEN_29;
  wire [1:0] GEN_30;
  reg [1:0] lastGrant;
  reg [31:0] GEN_41;
  wire [1:0] GEN_31;
  wire  T_823;
  wire  T_825;
  wire  T_827;
  wire  T_829;
  wire  T_830;
  wire  T_831;
  wire  T_834;
  wire  T_835;
  wire  T_836;
  wire  T_837;
  wire  T_838;
  wire  T_842;
  wire  T_844;
  wire  T_846;
  wire  T_848;
  wire  T_850;
  wire  T_852;
  wire  T_856;
  wire  T_857;
  wire  T_858;
  wire  T_859;
  wire  T_860;
  wire  T_862;
  wire  T_863;
  wire  T_864;
  wire  T_866;
  wire  T_867;
  wire  T_868;
  wire  T_870;
  wire  T_871;
  wire  T_872;
  wire  T_874;
  wire  T_875;
  wire  T_876;
  wire [1:0] GEN_32;
  wire [1:0] GEN_33;
  wire [1:0] GEN_34;
  wire [1:0] GEN_35;
  wire [1:0] GEN_36;
  wire [1:0] GEN_37;
  assign io_in_0_ready = T_864;
  assign io_in_1_ready = T_868;
  assign io_in_2_ready = T_872;
  assign io_in_3_ready = T_876;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_beat = GEN_1;
  assign io_out_bits_client_xact_id = GEN_2;
  assign io_out_bits_manager_xact_id = GEN_3;
  assign io_out_bits_is_builtin_type = GEN_4;
  assign io_out_bits_g_type = GEN_5;
  assign io_out_bits_data = GEN_6;
  assign io_chosen = GEN_30;
  assign choice = GEN_37;
  assign GEN_0 = GEN_9;
  assign GEN_7 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_8 = 2'h2 == io_chosen ? io_in_2_valid : GEN_7;
  assign GEN_9 = 2'h3 == io_chosen ? io_in_3_valid : GEN_8;
  assign GEN_1 = GEN_12;
  assign GEN_10 = 2'h1 == io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_11 = 2'h2 == io_chosen ? io_in_2_bits_addr_beat : GEN_10;
  assign GEN_12 = 2'h3 == io_chosen ? io_in_3_bits_addr_beat : GEN_11;
  assign GEN_2 = GEN_15;
  assign GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_14 = 2'h2 == io_chosen ? io_in_2_bits_client_xact_id : GEN_13;
  assign GEN_15 = 2'h3 == io_chosen ? io_in_3_bits_client_xact_id : GEN_14;
  assign GEN_3 = GEN_18;
  assign GEN_16 = 2'h1 == io_chosen ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign GEN_17 = 2'h2 == io_chosen ? io_in_2_bits_manager_xact_id : GEN_16;
  assign GEN_18 = 2'h3 == io_chosen ? io_in_3_bits_manager_xact_id : GEN_17;
  assign GEN_4 = GEN_21;
  assign GEN_19 = 2'h1 == io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_20 = 2'h2 == io_chosen ? io_in_2_bits_is_builtin_type : GEN_19;
  assign GEN_21 = 2'h3 == io_chosen ? io_in_3_bits_is_builtin_type : GEN_20;
  assign GEN_5 = GEN_24;
  assign GEN_22 = 2'h1 == io_chosen ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign GEN_23 = 2'h2 == io_chosen ? io_in_2_bits_g_type : GEN_22;
  assign GEN_24 = 2'h3 == io_chosen ? io_in_3_bits_g_type : GEN_23;
  assign GEN_6 = GEN_27;
  assign GEN_25 = 2'h1 == io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_26 = 2'h2 == io_chosen ? io_in_2_bits_data : GEN_25;
  assign GEN_27 = 2'h3 == io_chosen ? io_in_3_bits_data : GEN_26;
  assign T_798 = T_794 != 3'h0;
  assign T_806_0 = 3'h5;
  assign GEN_38 = {{1'd0}, T_806_0};
  assign T_808 = io_out_bits_g_type == GEN_38;
  assign T_809 = io_out_bits_g_type == 4'h0;
  assign T_810 = io_out_bits_is_builtin_type ? T_808 : T_809;
  assign T_812 = io_out_ready & io_out_valid;
  assign T_813 = T_812 & T_810;
  assign T_817 = T_794 + 3'h1;
  assign T_818 = T_817[2:0];
  assign GEN_28 = T_813 ? io_chosen : T_796;
  assign GEN_29 = T_813 ? T_818 : T_794;
  assign GEN_30 = T_798 ? T_796 : choice;
  assign GEN_31 = T_812 ? io_chosen : lastGrant;
  assign T_823 = 2'h1 > lastGrant;
  assign T_825 = 2'h2 > lastGrant;
  assign T_827 = 2'h3 > lastGrant;
  assign T_829 = io_in_1_valid & T_823;
  assign T_830 = io_in_2_valid & T_825;
  assign T_831 = io_in_3_valid & T_827;
  assign T_834 = T_829 | T_830;
  assign T_835 = T_834 | T_831;
  assign T_836 = T_835 | io_in_0_valid;
  assign T_837 = T_836 | io_in_1_valid;
  assign T_838 = T_837 | io_in_2_valid;
  assign T_842 = T_829 == 1'h0;
  assign T_844 = T_834 == 1'h0;
  assign T_846 = T_835 == 1'h0;
  assign T_848 = T_836 == 1'h0;
  assign T_850 = T_837 == 1'h0;
  assign T_852 = T_838 == 1'h0;
  assign T_856 = T_823 | T_848;
  assign T_857 = T_842 & T_825;
  assign T_858 = T_857 | T_850;
  assign T_859 = T_844 & T_827;
  assign T_860 = T_859 | T_852;
  assign T_862 = T_796 == 2'h0;
  assign T_863 = T_798 ? T_862 : T_846;
  assign T_864 = T_863 & io_out_ready;
  assign T_866 = T_796 == 2'h1;
  assign T_867 = T_798 ? T_866 : T_856;
  assign T_868 = T_867 & io_out_ready;
  assign T_870 = T_796 == 2'h2;
  assign T_871 = T_798 ? T_870 : T_858;
  assign T_872 = T_871 & io_out_ready;
  assign T_874 = T_796 == 2'h3;
  assign T_875 = T_798 ? T_874 : T_860;
  assign T_876 = T_875 & io_out_ready;
  assign GEN_32 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_33 = io_in_1_valid ? 2'h1 : GEN_32;
  assign GEN_34 = io_in_0_valid ? 2'h0 : GEN_33;
  assign GEN_35 = T_831 ? 2'h3 : GEN_34;
  assign GEN_36 = T_830 ? 2'h2 : GEN_35;
  assign GEN_37 = T_829 ? 2'h1 : GEN_36;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_39 = {1{$random}};
  T_794 = GEN_39[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_40 = {1{$random}};
  T_796 = GEN_40[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_41 = {1{$random}};
  lastGrant = GEN_41[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_794 <= 3'h0;
    end else begin
      if(T_813) begin
        T_794 <= T_818;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_813) begin
        T_796 <= io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_812) begin
        lastGrant <= io_chosen;
      end
    end
  end
endmodule
module ClientUncachedTileLinkIORouter_1(
  input   clk,
  input   reset,
  output  io_in_acquire_ready,
  input   io_in_acquire_valid,
  input  [25:0] io_in_acquire_bits_addr_block,
  input  [1:0] io_in_acquire_bits_client_xact_id,
  input  [2:0] io_in_acquire_bits_addr_beat,
  input   io_in_acquire_bits_is_builtin_type,
  input  [2:0] io_in_acquire_bits_a_type,
  input  [11:0] io_in_acquire_bits_union,
  input  [63:0] io_in_acquire_bits_data,
  input   io_in_grant_ready,
  output  io_in_grant_valid,
  output [2:0] io_in_grant_bits_addr_beat,
  output [1:0] io_in_grant_bits_client_xact_id,
  output  io_in_grant_bits_manager_xact_id,
  output  io_in_grant_bits_is_builtin_type,
  output [3:0] io_in_grant_bits_g_type,
  output [63:0] io_in_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [11:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [11:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data,
  input   io_out_2_acquire_ready,
  output  io_out_2_acquire_valid,
  output [25:0] io_out_2_acquire_bits_addr_block,
  output [1:0] io_out_2_acquire_bits_client_xact_id,
  output [2:0] io_out_2_acquire_bits_addr_beat,
  output  io_out_2_acquire_bits_is_builtin_type,
  output [2:0] io_out_2_acquire_bits_a_type,
  output [11:0] io_out_2_acquire_bits_union,
  output [63:0] io_out_2_acquire_bits_data,
  output  io_out_2_grant_ready,
  input   io_out_2_grant_valid,
  input  [2:0] io_out_2_grant_bits_addr_beat,
  input  [1:0] io_out_2_grant_bits_client_xact_id,
  input   io_out_2_grant_bits_manager_xact_id,
  input   io_out_2_grant_bits_is_builtin_type,
  input  [3:0] io_out_2_grant_bits_g_type,
  input  [63:0] io_out_2_grant_bits_data,
  input   io_out_3_acquire_ready,
  output  io_out_3_acquire_valid,
  output [25:0] io_out_3_acquire_bits_addr_block,
  output [1:0] io_out_3_acquire_bits_client_xact_id,
  output [2:0] io_out_3_acquire_bits_addr_beat,
  output  io_out_3_acquire_bits_is_builtin_type,
  output [2:0] io_out_3_acquire_bits_a_type,
  output [11:0] io_out_3_acquire_bits_union,
  output [63:0] io_out_3_acquire_bits_data,
  output  io_out_3_grant_ready,
  input   io_out_3_grant_valid,
  input  [2:0] io_out_3_grant_bits_addr_beat,
  input  [1:0] io_out_3_grant_bits_client_xact_id,
  input   io_out_3_grant_bits_manager_xact_id,
  input   io_out_3_grant_bits_is_builtin_type,
  input  [3:0] io_out_3_grant_bits_g_type,
  input  [63:0] io_out_3_grant_bits_data
);
  wire [2:0] T_1855_0;
  wire [2:0] T_1855_1;
  wire  T_1857;
  wire  T_1858;
  wire  T_1859;
  wire  T_1860;
  wire [2:0] T_1861;
  wire [2:0] T_1863;
  wire [28:0] T_1864;
  wire [31:0] T_1865;
  wire  T_1869;
  wire  T_1872;
  wire  T_1874;
  wire  T_1875;
  wire  T_1877;
  wire  T_1879;
  wire  T_1880;
  wire  T_1882;
  wire  T_1884;
  wire  T_1885;
  wire [1:0] T_1886;
  wire [1:0] T_1887;
  wire [3:0] acq_route;
  wire  T_1889;
  wire  T_1890;
  wire  GEN_0;
  wire  T_1892;
  wire  T_1893;
  wire  GEN_1;
  wire  T_1895;
  wire  T_1896;
  wire  GEN_2;
  wire  T_1898;
  wire  T_1899;
  wire  GEN_3;
  wire  gnt_arb_clk;
  wire  gnt_arb_reset;
  wire  gnt_arb_io_in_0_ready;
  wire  gnt_arb_io_in_0_valid;
  wire [2:0] gnt_arb_io_in_0_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_0_bits_client_xact_id;
  wire  gnt_arb_io_in_0_bits_manager_xact_id;
  wire  gnt_arb_io_in_0_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_0_bits_g_type;
  wire [63:0] gnt_arb_io_in_0_bits_data;
  wire  gnt_arb_io_in_1_ready;
  wire  gnt_arb_io_in_1_valid;
  wire [2:0] gnt_arb_io_in_1_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_1_bits_client_xact_id;
  wire  gnt_arb_io_in_1_bits_manager_xact_id;
  wire  gnt_arb_io_in_1_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_1_bits_g_type;
  wire [63:0] gnt_arb_io_in_1_bits_data;
  wire  gnt_arb_io_in_2_ready;
  wire  gnt_arb_io_in_2_valid;
  wire [2:0] gnt_arb_io_in_2_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_2_bits_client_xact_id;
  wire  gnt_arb_io_in_2_bits_manager_xact_id;
  wire  gnt_arb_io_in_2_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_2_bits_g_type;
  wire [63:0] gnt_arb_io_in_2_bits_data;
  wire  gnt_arb_io_in_3_ready;
  wire  gnt_arb_io_in_3_valid;
  wire [2:0] gnt_arb_io_in_3_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_3_bits_client_xact_id;
  wire  gnt_arb_io_in_3_bits_manager_xact_id;
  wire  gnt_arb_io_in_3_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_3_bits_g_type;
  wire [63:0] gnt_arb_io_in_3_bits_data;
  wire  gnt_arb_io_out_ready;
  wire  gnt_arb_io_out_valid;
  wire [2:0] gnt_arb_io_out_bits_addr_beat;
  wire [1:0] gnt_arb_io_out_bits_client_xact_id;
  wire  gnt_arb_io_out_bits_manager_xact_id;
  wire  gnt_arb_io_out_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_out_bits_g_type;
  wire [63:0] gnt_arb_io_out_bits_data;
  wire [1:0] gnt_arb_io_chosen;
  wire  T_1924;
  wire  T_1926;
  wire  T_1927;
  wire  T_1928;
  wire  T_1930;
  LockingRRArbiter_7 gnt_arb (
    .clk(gnt_arb_clk),
    .reset(gnt_arb_reset),
    .io_in_0_ready(gnt_arb_io_in_0_ready),
    .io_in_0_valid(gnt_arb_io_in_0_valid),
    .io_in_0_bits_addr_beat(gnt_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(gnt_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(gnt_arb_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(gnt_arb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(gnt_arb_io_in_0_bits_g_type),
    .io_in_0_bits_data(gnt_arb_io_in_0_bits_data),
    .io_in_1_ready(gnt_arb_io_in_1_ready),
    .io_in_1_valid(gnt_arb_io_in_1_valid),
    .io_in_1_bits_addr_beat(gnt_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_client_xact_id(gnt_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_manager_xact_id(gnt_arb_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_is_builtin_type(gnt_arb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_g_type(gnt_arb_io_in_1_bits_g_type),
    .io_in_1_bits_data(gnt_arb_io_in_1_bits_data),
    .io_in_2_ready(gnt_arb_io_in_2_ready),
    .io_in_2_valid(gnt_arb_io_in_2_valid),
    .io_in_2_bits_addr_beat(gnt_arb_io_in_2_bits_addr_beat),
    .io_in_2_bits_client_xact_id(gnt_arb_io_in_2_bits_client_xact_id),
    .io_in_2_bits_manager_xact_id(gnt_arb_io_in_2_bits_manager_xact_id),
    .io_in_2_bits_is_builtin_type(gnt_arb_io_in_2_bits_is_builtin_type),
    .io_in_2_bits_g_type(gnt_arb_io_in_2_bits_g_type),
    .io_in_2_bits_data(gnt_arb_io_in_2_bits_data),
    .io_in_3_ready(gnt_arb_io_in_3_ready),
    .io_in_3_valid(gnt_arb_io_in_3_valid),
    .io_in_3_bits_addr_beat(gnt_arb_io_in_3_bits_addr_beat),
    .io_in_3_bits_client_xact_id(gnt_arb_io_in_3_bits_client_xact_id),
    .io_in_3_bits_manager_xact_id(gnt_arb_io_in_3_bits_manager_xact_id),
    .io_in_3_bits_is_builtin_type(gnt_arb_io_in_3_bits_is_builtin_type),
    .io_in_3_bits_g_type(gnt_arb_io_in_3_bits_g_type),
    .io_in_3_bits_data(gnt_arb_io_in_3_bits_data),
    .io_out_ready(gnt_arb_io_out_ready),
    .io_out_valid(gnt_arb_io_out_valid),
    .io_out_bits_addr_beat(gnt_arb_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(gnt_arb_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(gnt_arb_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(gnt_arb_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(gnt_arb_io_out_bits_g_type),
    .io_out_bits_data(gnt_arb_io_out_bits_data),
    .io_chosen(gnt_arb_io_chosen)
  );
  assign io_in_acquire_ready = GEN_3;
  assign io_in_grant_valid = gnt_arb_io_out_valid;
  assign io_in_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_in_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_in_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_in_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_in_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_in_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_out_0_acquire_valid = T_1890;
  assign io_out_0_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_0_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_0_grant_ready = gnt_arb_io_in_0_ready;
  assign io_out_1_acquire_valid = T_1893;
  assign io_out_1_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_1_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_1_grant_ready = gnt_arb_io_in_1_ready;
  assign io_out_2_acquire_valid = T_1896;
  assign io_out_2_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_2_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_2_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_2_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_2_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_2_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_2_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_2_grant_ready = gnt_arb_io_in_2_ready;
  assign io_out_3_acquire_valid = T_1899;
  assign io_out_3_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_3_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_3_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_3_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_3_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_3_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_3_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_3_grant_ready = gnt_arb_io_in_3_ready;
  assign T_1855_0 = 3'h0;
  assign T_1855_1 = 3'h4;
  assign T_1857 = io_in_acquire_bits_a_type == T_1855_0;
  assign T_1858 = io_in_acquire_bits_a_type == T_1855_1;
  assign T_1859 = T_1857 | T_1858;
  assign T_1860 = io_in_acquire_bits_is_builtin_type & T_1859;
  assign T_1861 = io_in_acquire_bits_union[11:9];
  assign T_1863 = T_1860 ? T_1861 : 3'h0;
  assign T_1864 = {io_in_acquire_bits_addr_block,io_in_acquire_bits_addr_beat};
  assign T_1865 = {T_1864,T_1863};
  assign T_1869 = T_1865 < 32'h1000;
  assign T_1872 = 32'h1000 <= T_1865;
  assign T_1874 = T_1865 < 32'h2000;
  assign T_1875 = T_1872 & T_1874;
  assign T_1877 = 32'h40000000 <= T_1865;
  assign T_1879 = T_1865 < 32'h44000000;
  assign T_1880 = T_1877 & T_1879;
  assign T_1882 = 32'h44000000 <= T_1865;
  assign T_1884 = T_1865 < 32'h48000000;
  assign T_1885 = T_1882 & T_1884;
  assign T_1886 = {T_1875,T_1869};
  assign T_1887 = {T_1885,T_1880};
  assign acq_route = {T_1887,T_1886};
  assign T_1889 = acq_route[0];
  assign T_1890 = io_in_acquire_valid & T_1889;
  assign GEN_0 = T_1889 ? io_out_0_acquire_ready : 1'h0;
  assign T_1892 = acq_route[1];
  assign T_1893 = io_in_acquire_valid & T_1892;
  assign GEN_1 = T_1892 ? io_out_1_acquire_ready : GEN_0;
  assign T_1895 = acq_route[2];
  assign T_1896 = io_in_acquire_valid & T_1895;
  assign GEN_2 = T_1895 ? io_out_2_acquire_ready : GEN_1;
  assign T_1898 = acq_route[3];
  assign T_1899 = io_in_acquire_valid & T_1898;
  assign GEN_3 = T_1898 ? io_out_3_acquire_ready : GEN_2;
  assign gnt_arb_clk = clk;
  assign gnt_arb_reset = reset;
  assign gnt_arb_io_in_0_valid = io_out_0_grant_valid;
  assign gnt_arb_io_in_0_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign gnt_arb_io_in_0_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign gnt_arb_io_in_0_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_0_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_0_bits_g_type = io_out_0_grant_bits_g_type;
  assign gnt_arb_io_in_0_bits_data = io_out_0_grant_bits_data;
  assign gnt_arb_io_in_1_valid = io_out_1_grant_valid;
  assign gnt_arb_io_in_1_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign gnt_arb_io_in_1_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign gnt_arb_io_in_1_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_1_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_1_bits_g_type = io_out_1_grant_bits_g_type;
  assign gnt_arb_io_in_1_bits_data = io_out_1_grant_bits_data;
  assign gnt_arb_io_in_2_valid = io_out_2_grant_valid;
  assign gnt_arb_io_in_2_bits_addr_beat = io_out_2_grant_bits_addr_beat;
  assign gnt_arb_io_in_2_bits_client_xact_id = io_out_2_grant_bits_client_xact_id;
  assign gnt_arb_io_in_2_bits_manager_xact_id = io_out_2_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_2_bits_is_builtin_type = io_out_2_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_2_bits_g_type = io_out_2_grant_bits_g_type;
  assign gnt_arb_io_in_2_bits_data = io_out_2_grant_bits_data;
  assign gnt_arb_io_in_3_valid = io_out_3_grant_valid;
  assign gnt_arb_io_in_3_bits_addr_beat = io_out_3_grant_bits_addr_beat;
  assign gnt_arb_io_in_3_bits_client_xact_id = io_out_3_grant_bits_client_xact_id;
  assign gnt_arb_io_in_3_bits_manager_xact_id = io_out_3_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_3_bits_is_builtin_type = io_out_3_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_3_bits_g_type = io_out_3_grant_bits_g_type;
  assign gnt_arb_io_in_3_bits_data = io_out_3_grant_bits_data;
  assign gnt_arb_io_out_ready = io_in_grant_ready;
  assign T_1924 = io_in_acquire_valid == 1'h0;
  assign T_1926 = acq_route != 4'h0;
  assign T_1927 = T_1924 | T_1926;
  assign T_1928 = T_1927 | reset;
  assign T_1930 = T_1928 == 1'h0;
  always @(posedge clk) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1930) begin
          $fwrite(32'h80000002,"Assertion failed: No valid route\n    at Interconnect.scala:219 assert(!io.in.acquire.valid || acq_route.orR, ---No valid route---)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1930) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module ClientUncachedTileLinkIOCrossbar_1(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [11:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [11:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data,
  input   io_out_2_acquire_ready,
  output  io_out_2_acquire_valid,
  output [25:0] io_out_2_acquire_bits_addr_block,
  output [1:0] io_out_2_acquire_bits_client_xact_id,
  output [2:0] io_out_2_acquire_bits_addr_beat,
  output  io_out_2_acquire_bits_is_builtin_type,
  output [2:0] io_out_2_acquire_bits_a_type,
  output [11:0] io_out_2_acquire_bits_union,
  output [63:0] io_out_2_acquire_bits_data,
  output  io_out_2_grant_ready,
  input   io_out_2_grant_valid,
  input  [2:0] io_out_2_grant_bits_addr_beat,
  input  [1:0] io_out_2_grant_bits_client_xact_id,
  input   io_out_2_grant_bits_manager_xact_id,
  input   io_out_2_grant_bits_is_builtin_type,
  input  [3:0] io_out_2_grant_bits_g_type,
  input  [63:0] io_out_2_grant_bits_data,
  input   io_out_3_acquire_ready,
  output  io_out_3_acquire_valid,
  output [25:0] io_out_3_acquire_bits_addr_block,
  output [1:0] io_out_3_acquire_bits_client_xact_id,
  output [2:0] io_out_3_acquire_bits_addr_beat,
  output  io_out_3_acquire_bits_is_builtin_type,
  output [2:0] io_out_3_acquire_bits_a_type,
  output [11:0] io_out_3_acquire_bits_union,
  output [63:0] io_out_3_acquire_bits_data,
  output  io_out_3_grant_ready,
  input   io_out_3_grant_valid,
  input  [2:0] io_out_3_grant_bits_addr_beat,
  input  [1:0] io_out_3_grant_bits_client_xact_id,
  input   io_out_3_grant_bits_manager_xact_id,
  input   io_out_3_grant_bits_is_builtin_type,
  input  [3:0] io_out_3_grant_bits_g_type,
  input  [63:0] io_out_3_grant_bits_data
);
  wire  ClientUncachedTileLinkIORouter_1_1_clk;
  wire  ClientUncachedTileLinkIORouter_1_1_reset;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_ready;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_data;
  ClientUncachedTileLinkIORouter_1 ClientUncachedTileLinkIORouter_1_1 (
    .clk(ClientUncachedTileLinkIORouter_1_1_clk),
    .reset(ClientUncachedTileLinkIORouter_1_1_reset),
    .io_in_acquire_ready(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_ready),
    .io_in_acquire_valid(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_valid),
    .io_in_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_block),
    .io_in_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_client_xact_id),
    .io_in_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_beat),
    .io_in_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_is_builtin_type),
    .io_in_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_a_type),
    .io_in_acquire_bits_union(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_union),
    .io_in_acquire_bits_data(ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_data),
    .io_in_grant_ready(ClientUncachedTileLinkIORouter_1_1_io_in_grant_ready),
    .io_in_grant_valid(ClientUncachedTileLinkIORouter_1_1_io_in_grant_valid),
    .io_in_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_addr_beat),
    .io_in_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_client_xact_id),
    .io_in_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_manager_xact_id),
    .io_in_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_is_builtin_type),
    .io_in_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_g_type),
    .io_in_grant_bits_data(ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_data),
    .io_out_0_acquire_ready(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_ready),
    .io_out_0_grant_valid(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_ready),
    .io_out_1_grant_valid(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_data),
    .io_out_2_acquire_ready(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_ready),
    .io_out_2_acquire_valid(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_valid),
    .io_out_2_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_block),
    .io_out_2_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_client_xact_id),
    .io_out_2_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_beat),
    .io_out_2_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_is_builtin_type),
    .io_out_2_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_a_type),
    .io_out_2_acquire_bits_union(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_union),
    .io_out_2_acquire_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_data),
    .io_out_2_grant_ready(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_ready),
    .io_out_2_grant_valid(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_valid),
    .io_out_2_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_addr_beat),
    .io_out_2_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_client_xact_id),
    .io_out_2_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_manager_xact_id),
    .io_out_2_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_is_builtin_type),
    .io_out_2_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_g_type),
    .io_out_2_grant_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_data),
    .io_out_3_acquire_ready(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_ready),
    .io_out_3_acquire_valid(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_valid),
    .io_out_3_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_block),
    .io_out_3_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_client_xact_id),
    .io_out_3_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_beat),
    .io_out_3_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_is_builtin_type),
    .io_out_3_acquire_bits_a_type(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_a_type),
    .io_out_3_acquire_bits_union(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_union),
    .io_out_3_acquire_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_data),
    .io_out_3_grant_ready(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_ready),
    .io_out_3_grant_valid(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_valid),
    .io_out_3_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_addr_beat),
    .io_out_3_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_client_xact_id),
    .io_out_3_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_manager_xact_id),
    .io_out_3_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_is_builtin_type),
    .io_out_3_grant_bits_g_type(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_g_type),
    .io_out_3_grant_bits_data(ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_data)
  );
  assign io_in_0_acquire_ready = ClientUncachedTileLinkIORouter_1_1_io_in_acquire_ready;
  assign io_in_0_grant_valid = ClientUncachedTileLinkIORouter_1_1_io_in_grant_valid;
  assign io_in_0_grant_bits_addr_beat = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_g_type;
  assign io_in_0_grant_bits_data = ClientUncachedTileLinkIORouter_1_1_io_in_grant_bits_data;
  assign io_out_0_acquire_valid = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_union;
  assign io_out_0_acquire_bits_data = ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_bits_data;
  assign io_out_0_grant_ready = ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_ready;
  assign io_out_1_acquire_valid = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_valid;
  assign io_out_1_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_union;
  assign io_out_1_acquire_bits_data = ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_bits_data;
  assign io_out_1_grant_ready = ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_ready;
  assign io_out_2_acquire_valid = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_valid;
  assign io_out_2_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_block;
  assign io_out_2_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_client_xact_id;
  assign io_out_2_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_addr_beat;
  assign io_out_2_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_is_builtin_type;
  assign io_out_2_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_a_type;
  assign io_out_2_acquire_bits_union = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_union;
  assign io_out_2_acquire_bits_data = ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_bits_data;
  assign io_out_2_grant_ready = ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_ready;
  assign io_out_3_acquire_valid = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_valid;
  assign io_out_3_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_block;
  assign io_out_3_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_client_xact_id;
  assign io_out_3_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_addr_beat;
  assign io_out_3_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_is_builtin_type;
  assign io_out_3_acquire_bits_a_type = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_a_type;
  assign io_out_3_acquire_bits_union = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_union;
  assign io_out_3_acquire_bits_data = ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_bits_data;
  assign io_out_3_grant_ready = ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_ready;
  assign ClientUncachedTileLinkIORouter_1_1_clk = clk;
  assign ClientUncachedTileLinkIORouter_1_1_reset = reset;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_valid = io_in_0_acquire_valid;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_union = io_in_0_acquire_bits_union;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_acquire_bits_data = io_in_0_acquire_bits_data;
  assign ClientUncachedTileLinkIORouter_1_1_io_in_grant_ready = io_in_0_grant_ready;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_acquire_ready = io_out_0_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_valid = io_out_0_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_0_grant_bits_data = io_out_0_grant_bits_data;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_acquire_ready = io_out_1_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_valid = io_out_1_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_g_type = io_out_1_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_1_grant_bits_data = io_out_1_grant_bits_data;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_acquire_ready = io_out_2_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_valid = io_out_2_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_addr_beat = io_out_2_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_client_xact_id = io_out_2_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_manager_xact_id = io_out_2_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_is_builtin_type = io_out_2_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_g_type = io_out_2_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_2_grant_bits_data = io_out_2_grant_bits_data;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_acquire_ready = io_out_3_acquire_ready;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_valid = io_out_3_grant_valid;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_addr_beat = io_out_3_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_client_xact_id = io_out_3_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_manager_xact_id = io_out_3_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_is_builtin_type = io_out_3_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_g_type = io_out_3_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_1_1_io_out_3_grant_bits_data = io_out_3_grant_bits_data;
endmodule
module TileLinkRecursiveInterconnect_1(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [11:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [11:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data,
  input   io_out_2_acquire_ready,
  output  io_out_2_acquire_valid,
  output [25:0] io_out_2_acquire_bits_addr_block,
  output [1:0] io_out_2_acquire_bits_client_xact_id,
  output [2:0] io_out_2_acquire_bits_addr_beat,
  output  io_out_2_acquire_bits_is_builtin_type,
  output [2:0] io_out_2_acquire_bits_a_type,
  output [11:0] io_out_2_acquire_bits_union,
  output [63:0] io_out_2_acquire_bits_data,
  output  io_out_2_grant_ready,
  input   io_out_2_grant_valid,
  input  [2:0] io_out_2_grant_bits_addr_beat,
  input  [1:0] io_out_2_grant_bits_client_xact_id,
  input   io_out_2_grant_bits_manager_xact_id,
  input   io_out_2_grant_bits_is_builtin_type,
  input  [3:0] io_out_2_grant_bits_g_type,
  input  [63:0] io_out_2_grant_bits_data,
  input   io_out_3_acquire_ready,
  output  io_out_3_acquire_valid,
  output [25:0] io_out_3_acquire_bits_addr_block,
  output [1:0] io_out_3_acquire_bits_client_xact_id,
  output [2:0] io_out_3_acquire_bits_addr_beat,
  output  io_out_3_acquire_bits_is_builtin_type,
  output [2:0] io_out_3_acquire_bits_a_type,
  output [11:0] io_out_3_acquire_bits_union,
  output [63:0] io_out_3_acquire_bits_data,
  output  io_out_3_grant_ready,
  input   io_out_3_grant_valid,
  input  [2:0] io_out_3_grant_bits_addr_beat,
  input  [1:0] io_out_3_grant_bits_client_xact_id,
  input   io_out_3_grant_bits_manager_xact_id,
  input   io_out_3_grant_bits_is_builtin_type,
  input  [3:0] io_out_3_grant_bits_g_type,
  input  [63:0] io_out_3_grant_bits_data
);
  wire  xbar_clk;
  wire  xbar_reset;
  wire  xbar_io_in_0_acquire_ready;
  wire  xbar_io_in_0_acquire_valid;
  wire [25:0] xbar_io_in_0_acquire_bits_addr_block;
  wire [1:0] xbar_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_in_0_acquire_bits_addr_beat;
  wire  xbar_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_in_0_acquire_bits_a_type;
  wire [11:0] xbar_io_in_0_acquire_bits_union;
  wire [63:0] xbar_io_in_0_acquire_bits_data;
  wire  xbar_io_in_0_grant_ready;
  wire  xbar_io_in_0_grant_valid;
  wire [2:0] xbar_io_in_0_grant_bits_addr_beat;
  wire [1:0] xbar_io_in_0_grant_bits_client_xact_id;
  wire  xbar_io_in_0_grant_bits_manager_xact_id;
  wire  xbar_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_in_0_grant_bits_g_type;
  wire [63:0] xbar_io_in_0_grant_bits_data;
  wire  xbar_io_out_0_acquire_ready;
  wire  xbar_io_out_0_acquire_valid;
  wire [25:0] xbar_io_out_0_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_0_acquire_bits_addr_beat;
  wire  xbar_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_0_acquire_bits_a_type;
  wire [11:0] xbar_io_out_0_acquire_bits_union;
  wire [63:0] xbar_io_out_0_acquire_bits_data;
  wire  xbar_io_out_0_grant_ready;
  wire  xbar_io_out_0_grant_valid;
  wire [2:0] xbar_io_out_0_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_0_grant_bits_client_xact_id;
  wire  xbar_io_out_0_grant_bits_manager_xact_id;
  wire  xbar_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_0_grant_bits_g_type;
  wire [63:0] xbar_io_out_0_grant_bits_data;
  wire  xbar_io_out_1_acquire_ready;
  wire  xbar_io_out_1_acquire_valid;
  wire [25:0] xbar_io_out_1_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_1_acquire_bits_addr_beat;
  wire  xbar_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_1_acquire_bits_a_type;
  wire [11:0] xbar_io_out_1_acquire_bits_union;
  wire [63:0] xbar_io_out_1_acquire_bits_data;
  wire  xbar_io_out_1_grant_ready;
  wire  xbar_io_out_1_grant_valid;
  wire [2:0] xbar_io_out_1_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_1_grant_bits_client_xact_id;
  wire  xbar_io_out_1_grant_bits_manager_xact_id;
  wire  xbar_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_1_grant_bits_g_type;
  wire [63:0] xbar_io_out_1_grant_bits_data;
  wire  xbar_io_out_2_acquire_ready;
  wire  xbar_io_out_2_acquire_valid;
  wire [25:0] xbar_io_out_2_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_2_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_2_acquire_bits_addr_beat;
  wire  xbar_io_out_2_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_2_acquire_bits_a_type;
  wire [11:0] xbar_io_out_2_acquire_bits_union;
  wire [63:0] xbar_io_out_2_acquire_bits_data;
  wire  xbar_io_out_2_grant_ready;
  wire  xbar_io_out_2_grant_valid;
  wire [2:0] xbar_io_out_2_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_2_grant_bits_client_xact_id;
  wire  xbar_io_out_2_grant_bits_manager_xact_id;
  wire  xbar_io_out_2_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_2_grant_bits_g_type;
  wire [63:0] xbar_io_out_2_grant_bits_data;
  wire  xbar_io_out_3_acquire_ready;
  wire  xbar_io_out_3_acquire_valid;
  wire [25:0] xbar_io_out_3_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_3_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_3_acquire_bits_addr_beat;
  wire  xbar_io_out_3_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_3_acquire_bits_a_type;
  wire [11:0] xbar_io_out_3_acquire_bits_union;
  wire [63:0] xbar_io_out_3_acquire_bits_data;
  wire  xbar_io_out_3_grant_ready;
  wire  xbar_io_out_3_grant_valid;
  wire [2:0] xbar_io_out_3_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_3_grant_bits_client_xact_id;
  wire  xbar_io_out_3_grant_bits_manager_xact_id;
  wire  xbar_io_out_3_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_3_grant_bits_g_type;
  wire [63:0] xbar_io_out_3_grant_bits_data;
  ClientUncachedTileLinkIOCrossbar_1 xbar (
    .clk(xbar_clk),
    .reset(xbar_reset),
    .io_in_0_acquire_ready(xbar_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(xbar_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(xbar_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(xbar_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(xbar_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(xbar_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(xbar_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(xbar_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(xbar_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(xbar_io_in_0_grant_ready),
    .io_in_0_grant_valid(xbar_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(xbar_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(xbar_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(xbar_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(xbar_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(xbar_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(xbar_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(xbar_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(xbar_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(xbar_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(xbar_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(xbar_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(xbar_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(xbar_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(xbar_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(xbar_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(xbar_io_out_0_grant_ready),
    .io_out_0_grant_valid(xbar_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(xbar_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(xbar_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(xbar_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(xbar_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(xbar_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(xbar_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(xbar_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(xbar_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(xbar_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(xbar_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(xbar_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(xbar_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(xbar_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(xbar_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(xbar_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(xbar_io_out_1_grant_ready),
    .io_out_1_grant_valid(xbar_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(xbar_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(xbar_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(xbar_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(xbar_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(xbar_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(xbar_io_out_1_grant_bits_data),
    .io_out_2_acquire_ready(xbar_io_out_2_acquire_ready),
    .io_out_2_acquire_valid(xbar_io_out_2_acquire_valid),
    .io_out_2_acquire_bits_addr_block(xbar_io_out_2_acquire_bits_addr_block),
    .io_out_2_acquire_bits_client_xact_id(xbar_io_out_2_acquire_bits_client_xact_id),
    .io_out_2_acquire_bits_addr_beat(xbar_io_out_2_acquire_bits_addr_beat),
    .io_out_2_acquire_bits_is_builtin_type(xbar_io_out_2_acquire_bits_is_builtin_type),
    .io_out_2_acquire_bits_a_type(xbar_io_out_2_acquire_bits_a_type),
    .io_out_2_acquire_bits_union(xbar_io_out_2_acquire_bits_union),
    .io_out_2_acquire_bits_data(xbar_io_out_2_acquire_bits_data),
    .io_out_2_grant_ready(xbar_io_out_2_grant_ready),
    .io_out_2_grant_valid(xbar_io_out_2_grant_valid),
    .io_out_2_grant_bits_addr_beat(xbar_io_out_2_grant_bits_addr_beat),
    .io_out_2_grant_bits_client_xact_id(xbar_io_out_2_grant_bits_client_xact_id),
    .io_out_2_grant_bits_manager_xact_id(xbar_io_out_2_grant_bits_manager_xact_id),
    .io_out_2_grant_bits_is_builtin_type(xbar_io_out_2_grant_bits_is_builtin_type),
    .io_out_2_grant_bits_g_type(xbar_io_out_2_grant_bits_g_type),
    .io_out_2_grant_bits_data(xbar_io_out_2_grant_bits_data),
    .io_out_3_acquire_ready(xbar_io_out_3_acquire_ready),
    .io_out_3_acquire_valid(xbar_io_out_3_acquire_valid),
    .io_out_3_acquire_bits_addr_block(xbar_io_out_3_acquire_bits_addr_block),
    .io_out_3_acquire_bits_client_xact_id(xbar_io_out_3_acquire_bits_client_xact_id),
    .io_out_3_acquire_bits_addr_beat(xbar_io_out_3_acquire_bits_addr_beat),
    .io_out_3_acquire_bits_is_builtin_type(xbar_io_out_3_acquire_bits_is_builtin_type),
    .io_out_3_acquire_bits_a_type(xbar_io_out_3_acquire_bits_a_type),
    .io_out_3_acquire_bits_union(xbar_io_out_3_acquire_bits_union),
    .io_out_3_acquire_bits_data(xbar_io_out_3_acquire_bits_data),
    .io_out_3_grant_ready(xbar_io_out_3_grant_ready),
    .io_out_3_grant_valid(xbar_io_out_3_grant_valid),
    .io_out_3_grant_bits_addr_beat(xbar_io_out_3_grant_bits_addr_beat),
    .io_out_3_grant_bits_client_xact_id(xbar_io_out_3_grant_bits_client_xact_id),
    .io_out_3_grant_bits_manager_xact_id(xbar_io_out_3_grant_bits_manager_xact_id),
    .io_out_3_grant_bits_is_builtin_type(xbar_io_out_3_grant_bits_is_builtin_type),
    .io_out_3_grant_bits_g_type(xbar_io_out_3_grant_bits_g_type),
    .io_out_3_grant_bits_data(xbar_io_out_3_grant_bits_data)
  );
  assign io_in_0_acquire_ready = xbar_io_in_0_acquire_ready;
  assign io_in_0_grant_valid = xbar_io_in_0_grant_valid;
  assign io_in_0_grant_bits_addr_beat = xbar_io_in_0_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = xbar_io_in_0_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = xbar_io_in_0_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = xbar_io_in_0_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = xbar_io_in_0_grant_bits_g_type;
  assign io_in_0_grant_bits_data = xbar_io_in_0_grant_bits_data;
  assign io_out_0_acquire_valid = xbar_io_out_0_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = xbar_io_out_0_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = xbar_io_out_0_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = xbar_io_out_0_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = xbar_io_out_0_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = xbar_io_out_0_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = xbar_io_out_0_acquire_bits_union;
  assign io_out_0_acquire_bits_data = xbar_io_out_0_acquire_bits_data;
  assign io_out_0_grant_ready = xbar_io_out_0_grant_ready;
  assign io_out_1_acquire_valid = xbar_io_out_1_acquire_valid;
  assign io_out_1_acquire_bits_addr_block = xbar_io_out_1_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = xbar_io_out_1_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = xbar_io_out_1_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = xbar_io_out_1_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = xbar_io_out_1_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = xbar_io_out_1_acquire_bits_union;
  assign io_out_1_acquire_bits_data = xbar_io_out_1_acquire_bits_data;
  assign io_out_1_grant_ready = xbar_io_out_1_grant_ready;
  assign io_out_2_acquire_valid = xbar_io_out_2_acquire_valid;
  assign io_out_2_acquire_bits_addr_block = xbar_io_out_2_acquire_bits_addr_block;
  assign io_out_2_acquire_bits_client_xact_id = xbar_io_out_2_acquire_bits_client_xact_id;
  assign io_out_2_acquire_bits_addr_beat = xbar_io_out_2_acquire_bits_addr_beat;
  assign io_out_2_acquire_bits_is_builtin_type = xbar_io_out_2_acquire_bits_is_builtin_type;
  assign io_out_2_acquire_bits_a_type = xbar_io_out_2_acquire_bits_a_type;
  assign io_out_2_acquire_bits_union = xbar_io_out_2_acquire_bits_union;
  assign io_out_2_acquire_bits_data = xbar_io_out_2_acquire_bits_data;
  assign io_out_2_grant_ready = xbar_io_out_2_grant_ready;
  assign io_out_3_acquire_valid = xbar_io_out_3_acquire_valid;
  assign io_out_3_acquire_bits_addr_block = xbar_io_out_3_acquire_bits_addr_block;
  assign io_out_3_acquire_bits_client_xact_id = xbar_io_out_3_acquire_bits_client_xact_id;
  assign io_out_3_acquire_bits_addr_beat = xbar_io_out_3_acquire_bits_addr_beat;
  assign io_out_3_acquire_bits_is_builtin_type = xbar_io_out_3_acquire_bits_is_builtin_type;
  assign io_out_3_acquire_bits_a_type = xbar_io_out_3_acquire_bits_a_type;
  assign io_out_3_acquire_bits_union = xbar_io_out_3_acquire_bits_union;
  assign io_out_3_acquire_bits_data = xbar_io_out_3_acquire_bits_data;
  assign io_out_3_grant_ready = xbar_io_out_3_grant_ready;
  assign xbar_clk = clk;
  assign xbar_reset = reset;
  assign xbar_io_in_0_acquire_valid = io_in_0_acquire_valid;
  assign xbar_io_in_0_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign xbar_io_in_0_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign xbar_io_in_0_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign xbar_io_in_0_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign xbar_io_in_0_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign xbar_io_in_0_acquire_bits_union = io_in_0_acquire_bits_union;
  assign xbar_io_in_0_acquire_bits_data = io_in_0_acquire_bits_data;
  assign xbar_io_in_0_grant_ready = io_in_0_grant_ready;
  assign xbar_io_out_0_acquire_ready = io_out_0_acquire_ready;
  assign xbar_io_out_0_grant_valid = io_out_0_grant_valid;
  assign xbar_io_out_0_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign xbar_io_out_0_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign xbar_io_out_0_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign xbar_io_out_0_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign xbar_io_out_0_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign xbar_io_out_0_grant_bits_data = io_out_0_grant_bits_data;
  assign xbar_io_out_1_acquire_ready = io_out_1_acquire_ready;
  assign xbar_io_out_1_grant_valid = io_out_1_grant_valid;
  assign xbar_io_out_1_grant_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign xbar_io_out_1_grant_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign xbar_io_out_1_grant_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign xbar_io_out_1_grant_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign xbar_io_out_1_grant_bits_g_type = io_out_1_grant_bits_g_type;
  assign xbar_io_out_1_grant_bits_data = io_out_1_grant_bits_data;
  assign xbar_io_out_2_acquire_ready = io_out_2_acquire_ready;
  assign xbar_io_out_2_grant_valid = io_out_2_grant_valid;
  assign xbar_io_out_2_grant_bits_addr_beat = io_out_2_grant_bits_addr_beat;
  assign xbar_io_out_2_grant_bits_client_xact_id = io_out_2_grant_bits_client_xact_id;
  assign xbar_io_out_2_grant_bits_manager_xact_id = io_out_2_grant_bits_manager_xact_id;
  assign xbar_io_out_2_grant_bits_is_builtin_type = io_out_2_grant_bits_is_builtin_type;
  assign xbar_io_out_2_grant_bits_g_type = io_out_2_grant_bits_g_type;
  assign xbar_io_out_2_grant_bits_data = io_out_2_grant_bits_data;
  assign xbar_io_out_3_acquire_ready = io_out_3_acquire_ready;
  assign xbar_io_out_3_grant_valid = io_out_3_grant_valid;
  assign xbar_io_out_3_grant_bits_addr_beat = io_out_3_grant_bits_addr_beat;
  assign xbar_io_out_3_grant_bits_client_xact_id = io_out_3_grant_bits_client_xact_id;
  assign xbar_io_out_3_grant_bits_manager_xact_id = io_out_3_grant_bits_manager_xact_id;
  assign xbar_io_out_3_grant_bits_is_builtin_type = io_out_3_grant_bits_is_builtin_type;
  assign xbar_io_out_3_grant_bits_g_type = io_out_3_grant_bits_g_type;
  assign xbar_io_out_3_grant_bits_data = io_out_3_grant_bits_data;
endmodule
module TileLinkRecursiveInterconnect(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [11:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [11:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data,
  input   io_out_2_acquire_ready,
  output  io_out_2_acquire_valid,
  output [25:0] io_out_2_acquire_bits_addr_block,
  output [1:0] io_out_2_acquire_bits_client_xact_id,
  output [2:0] io_out_2_acquire_bits_addr_beat,
  output  io_out_2_acquire_bits_is_builtin_type,
  output [2:0] io_out_2_acquire_bits_a_type,
  output [11:0] io_out_2_acquire_bits_union,
  output [63:0] io_out_2_acquire_bits_data,
  output  io_out_2_grant_ready,
  input   io_out_2_grant_valid,
  input  [2:0] io_out_2_grant_bits_addr_beat,
  input  [1:0] io_out_2_grant_bits_client_xact_id,
  input   io_out_2_grant_bits_manager_xact_id,
  input   io_out_2_grant_bits_is_builtin_type,
  input  [3:0] io_out_2_grant_bits_g_type,
  input  [63:0] io_out_2_grant_bits_data,
  input   io_out_3_acquire_ready,
  output  io_out_3_acquire_valid,
  output [25:0] io_out_3_acquire_bits_addr_block,
  output [1:0] io_out_3_acquire_bits_client_xact_id,
  output [2:0] io_out_3_acquire_bits_addr_beat,
  output  io_out_3_acquire_bits_is_builtin_type,
  output [2:0] io_out_3_acquire_bits_a_type,
  output [11:0] io_out_3_acquire_bits_union,
  output [63:0] io_out_3_acquire_bits_data,
  output  io_out_3_grant_ready,
  input   io_out_3_grant_valid,
  input  [2:0] io_out_3_grant_bits_addr_beat,
  input  [1:0] io_out_3_grant_bits_client_xact_id,
  input   io_out_3_grant_bits_manager_xact_id,
  input   io_out_3_grant_bits_is_builtin_type,
  input  [3:0] io_out_3_grant_bits_g_type,
  input  [63:0] io_out_3_grant_bits_data,
  input   io_out_4_acquire_ready,
  output  io_out_4_acquire_valid,
  output [25:0] io_out_4_acquire_bits_addr_block,
  output [1:0] io_out_4_acquire_bits_client_xact_id,
  output [2:0] io_out_4_acquire_bits_addr_beat,
  output  io_out_4_acquire_bits_is_builtin_type,
  output [2:0] io_out_4_acquire_bits_a_type,
  output [11:0] io_out_4_acquire_bits_union,
  output [63:0] io_out_4_acquire_bits_data,
  output  io_out_4_grant_ready,
  input   io_out_4_grant_valid,
  input  [2:0] io_out_4_grant_bits_addr_beat,
  input  [1:0] io_out_4_grant_bits_client_xact_id,
  input   io_out_4_grant_bits_manager_xact_id,
  input   io_out_4_grant_bits_is_builtin_type,
  input  [3:0] io_out_4_grant_bits_g_type,
  input  [63:0] io_out_4_grant_bits_data
);
  wire  xbar_clk;
  wire  xbar_reset;
  wire  xbar_io_in_0_acquire_ready;
  wire  xbar_io_in_0_acquire_valid;
  wire [25:0] xbar_io_in_0_acquire_bits_addr_block;
  wire [1:0] xbar_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_in_0_acquire_bits_addr_beat;
  wire  xbar_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_in_0_acquire_bits_a_type;
  wire [11:0] xbar_io_in_0_acquire_bits_union;
  wire [63:0] xbar_io_in_0_acquire_bits_data;
  wire  xbar_io_in_0_grant_ready;
  wire  xbar_io_in_0_grant_valid;
  wire [2:0] xbar_io_in_0_grant_bits_addr_beat;
  wire [1:0] xbar_io_in_0_grant_bits_client_xact_id;
  wire  xbar_io_in_0_grant_bits_manager_xact_id;
  wire  xbar_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_in_0_grant_bits_g_type;
  wire [63:0] xbar_io_in_0_grant_bits_data;
  wire  xbar_io_out_0_acquire_ready;
  wire  xbar_io_out_0_acquire_valid;
  wire [25:0] xbar_io_out_0_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_0_acquire_bits_addr_beat;
  wire  xbar_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_0_acquire_bits_a_type;
  wire [11:0] xbar_io_out_0_acquire_bits_union;
  wire [63:0] xbar_io_out_0_acquire_bits_data;
  wire  xbar_io_out_0_grant_ready;
  wire  xbar_io_out_0_grant_valid;
  wire [2:0] xbar_io_out_0_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_0_grant_bits_client_xact_id;
  wire  xbar_io_out_0_grant_bits_manager_xact_id;
  wire  xbar_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_0_grant_bits_g_type;
  wire [63:0] xbar_io_out_0_grant_bits_data;
  wire  xbar_io_out_1_acquire_ready;
  wire  xbar_io_out_1_acquire_valid;
  wire [25:0] xbar_io_out_1_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_1_acquire_bits_addr_beat;
  wire  xbar_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_1_acquire_bits_a_type;
  wire [11:0] xbar_io_out_1_acquire_bits_union;
  wire [63:0] xbar_io_out_1_acquire_bits_data;
  wire  xbar_io_out_1_grant_ready;
  wire  xbar_io_out_1_grant_valid;
  wire [2:0] xbar_io_out_1_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_1_grant_bits_client_xact_id;
  wire  xbar_io_out_1_grant_bits_manager_xact_id;
  wire  xbar_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_1_grant_bits_g_type;
  wire [63:0] xbar_io_out_1_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_clk;
  wire  TileLinkRecursiveInterconnect_1_1_reset;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_grant_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_grant_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_grant_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_grant_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_grant_ready;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_data;
  ClientUncachedTileLinkIOCrossbar xbar (
    .clk(xbar_clk),
    .reset(xbar_reset),
    .io_in_0_acquire_ready(xbar_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(xbar_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(xbar_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(xbar_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(xbar_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(xbar_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(xbar_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(xbar_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(xbar_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(xbar_io_in_0_grant_ready),
    .io_in_0_grant_valid(xbar_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(xbar_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(xbar_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(xbar_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(xbar_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(xbar_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(xbar_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(xbar_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(xbar_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(xbar_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(xbar_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(xbar_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(xbar_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(xbar_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(xbar_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(xbar_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(xbar_io_out_0_grant_ready),
    .io_out_0_grant_valid(xbar_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(xbar_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(xbar_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(xbar_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(xbar_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(xbar_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(xbar_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(xbar_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(xbar_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(xbar_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(xbar_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(xbar_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(xbar_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(xbar_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(xbar_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(xbar_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(xbar_io_out_1_grant_ready),
    .io_out_1_grant_valid(xbar_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(xbar_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(xbar_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(xbar_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(xbar_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(xbar_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(xbar_io_out_1_grant_bits_data)
  );
  TileLinkRecursiveInterconnect_1 TileLinkRecursiveInterconnect_1_1 (
    .clk(TileLinkRecursiveInterconnect_1_1_clk),
    .reset(TileLinkRecursiveInterconnect_1_1_reset),
    .io_in_0_acquire_ready(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_ready),
    .io_in_0_grant_valid(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_ready),
    .io_out_0_grant_valid(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_ready),
    .io_out_1_grant_valid(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_data),
    .io_out_2_acquire_ready(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_ready),
    .io_out_2_acquire_valid(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_valid),
    .io_out_2_acquire_bits_addr_block(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_block),
    .io_out_2_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_client_xact_id),
    .io_out_2_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_beat),
    .io_out_2_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_is_builtin_type),
    .io_out_2_acquire_bits_a_type(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_a_type),
    .io_out_2_acquire_bits_union(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_union),
    .io_out_2_acquire_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_data),
    .io_out_2_grant_ready(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_ready),
    .io_out_2_grant_valid(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_valid),
    .io_out_2_grant_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_addr_beat),
    .io_out_2_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_client_xact_id),
    .io_out_2_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_manager_xact_id),
    .io_out_2_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_is_builtin_type),
    .io_out_2_grant_bits_g_type(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_g_type),
    .io_out_2_grant_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_data),
    .io_out_3_acquire_ready(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_ready),
    .io_out_3_acquire_valid(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_valid),
    .io_out_3_acquire_bits_addr_block(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_block),
    .io_out_3_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_client_xact_id),
    .io_out_3_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_beat),
    .io_out_3_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_is_builtin_type),
    .io_out_3_acquire_bits_a_type(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_a_type),
    .io_out_3_acquire_bits_union(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_union),
    .io_out_3_acquire_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_data),
    .io_out_3_grant_ready(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_ready),
    .io_out_3_grant_valid(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_valid),
    .io_out_3_grant_bits_addr_beat(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_addr_beat),
    .io_out_3_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_client_xact_id),
    .io_out_3_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_manager_xact_id),
    .io_out_3_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_is_builtin_type),
    .io_out_3_grant_bits_g_type(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_g_type),
    .io_out_3_grant_bits_data(TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_data)
  );
  assign io_in_0_acquire_ready = xbar_io_in_0_acquire_ready;
  assign io_in_0_grant_valid = xbar_io_in_0_grant_valid;
  assign io_in_0_grant_bits_addr_beat = xbar_io_in_0_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = xbar_io_in_0_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = xbar_io_in_0_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = xbar_io_in_0_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = xbar_io_in_0_grant_bits_g_type;
  assign io_in_0_grant_bits_data = xbar_io_in_0_grant_bits_data;
  assign io_out_0_acquire_valid = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_union;
  assign io_out_0_acquire_bits_data = TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_bits_data;
  assign io_out_0_grant_ready = TileLinkRecursiveInterconnect_1_1_io_out_0_grant_ready;
  assign io_out_1_acquire_valid = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_valid;
  assign io_out_1_acquire_bits_addr_block = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_union;
  assign io_out_1_acquire_bits_data = TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_bits_data;
  assign io_out_1_grant_ready = TileLinkRecursiveInterconnect_1_1_io_out_1_grant_ready;
  assign io_out_2_acquire_valid = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_valid;
  assign io_out_2_acquire_bits_addr_block = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_block;
  assign io_out_2_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_client_xact_id;
  assign io_out_2_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_addr_beat;
  assign io_out_2_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_is_builtin_type;
  assign io_out_2_acquire_bits_a_type = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_a_type;
  assign io_out_2_acquire_bits_union = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_union;
  assign io_out_2_acquire_bits_data = TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_bits_data;
  assign io_out_2_grant_ready = TileLinkRecursiveInterconnect_1_1_io_out_2_grant_ready;
  assign io_out_3_acquire_valid = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_valid;
  assign io_out_3_acquire_bits_addr_block = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_block;
  assign io_out_3_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_client_xact_id;
  assign io_out_3_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_addr_beat;
  assign io_out_3_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_is_builtin_type;
  assign io_out_3_acquire_bits_a_type = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_a_type;
  assign io_out_3_acquire_bits_union = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_union;
  assign io_out_3_acquire_bits_data = TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_bits_data;
  assign io_out_3_grant_ready = TileLinkRecursiveInterconnect_1_1_io_out_3_grant_ready;
  assign io_out_4_acquire_valid = xbar_io_out_1_acquire_valid;
  assign io_out_4_acquire_bits_addr_block = xbar_io_out_1_acquire_bits_addr_block;
  assign io_out_4_acquire_bits_client_xact_id = xbar_io_out_1_acquire_bits_client_xact_id;
  assign io_out_4_acquire_bits_addr_beat = xbar_io_out_1_acquire_bits_addr_beat;
  assign io_out_4_acquire_bits_is_builtin_type = xbar_io_out_1_acquire_bits_is_builtin_type;
  assign io_out_4_acquire_bits_a_type = xbar_io_out_1_acquire_bits_a_type;
  assign io_out_4_acquire_bits_union = xbar_io_out_1_acquire_bits_union;
  assign io_out_4_acquire_bits_data = xbar_io_out_1_acquire_bits_data;
  assign io_out_4_grant_ready = xbar_io_out_1_grant_ready;
  assign xbar_clk = clk;
  assign xbar_reset = reset;
  assign xbar_io_in_0_acquire_valid = io_in_0_acquire_valid;
  assign xbar_io_in_0_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign xbar_io_in_0_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign xbar_io_in_0_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign xbar_io_in_0_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign xbar_io_in_0_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign xbar_io_in_0_acquire_bits_union = io_in_0_acquire_bits_union;
  assign xbar_io_in_0_acquire_bits_data = io_in_0_acquire_bits_data;
  assign xbar_io_in_0_grant_ready = io_in_0_grant_ready;
  assign xbar_io_out_0_acquire_ready = TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_ready;
  assign xbar_io_out_0_grant_valid = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_valid;
  assign xbar_io_out_0_grant_bits_addr_beat = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_addr_beat;
  assign xbar_io_out_0_grant_bits_client_xact_id = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_client_xact_id;
  assign xbar_io_out_0_grant_bits_manager_xact_id = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_manager_xact_id;
  assign xbar_io_out_0_grant_bits_is_builtin_type = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_is_builtin_type;
  assign xbar_io_out_0_grant_bits_g_type = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_g_type;
  assign xbar_io_out_0_grant_bits_data = TileLinkRecursiveInterconnect_1_1_io_in_0_grant_bits_data;
  assign xbar_io_out_1_acquire_ready = io_out_4_acquire_ready;
  assign xbar_io_out_1_grant_valid = io_out_4_grant_valid;
  assign xbar_io_out_1_grant_bits_addr_beat = io_out_4_grant_bits_addr_beat;
  assign xbar_io_out_1_grant_bits_client_xact_id = io_out_4_grant_bits_client_xact_id;
  assign xbar_io_out_1_grant_bits_manager_xact_id = io_out_4_grant_bits_manager_xact_id;
  assign xbar_io_out_1_grant_bits_is_builtin_type = io_out_4_grant_bits_is_builtin_type;
  assign xbar_io_out_1_grant_bits_g_type = io_out_4_grant_bits_g_type;
  assign xbar_io_out_1_grant_bits_data = io_out_4_grant_bits_data;
  assign TileLinkRecursiveInterconnect_1_1_clk = clk;
  assign TileLinkRecursiveInterconnect_1_1_reset = reset;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_valid = xbar_io_out_0_acquire_valid;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_block = xbar_io_out_0_acquire_bits_addr_block;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_client_xact_id = xbar_io_out_0_acquire_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_addr_beat = xbar_io_out_0_acquire_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_is_builtin_type = xbar_io_out_0_acquire_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_a_type = xbar_io_out_0_acquire_bits_a_type;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_union = xbar_io_out_0_acquire_bits_union;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_acquire_bits_data = xbar_io_out_0_acquire_bits_data;
  assign TileLinkRecursiveInterconnect_1_1_io_in_0_grant_ready = xbar_io_out_0_grant_ready;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_acquire_ready = io_out_0_acquire_ready;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_valid = io_out_0_grant_valid;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_0_grant_bits_data = io_out_0_grant_bits_data;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_acquire_ready = io_out_1_acquire_ready;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_valid = io_out_1_grant_valid;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_g_type = io_out_1_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_1_grant_bits_data = io_out_1_grant_bits_data;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_acquire_ready = io_out_2_acquire_ready;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_valid = io_out_2_grant_valid;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_addr_beat = io_out_2_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_client_xact_id = io_out_2_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_manager_xact_id = io_out_2_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_is_builtin_type = io_out_2_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_g_type = io_out_2_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_2_grant_bits_data = io_out_2_grant_bits_data;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_acquire_ready = io_out_3_acquire_ready;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_valid = io_out_3_grant_valid;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_addr_beat = io_out_3_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_client_xact_id = io_out_3_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_manager_xact_id = io_out_3_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_is_builtin_type = io_out_3_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_g_type = io_out_3_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_1_1_io_out_3_grant_bits_data = io_out_3_grant_bits_data;
endmodule
module PLIC(
  input   clk,
  input   reset,
  input   io_devices_0_valid,
  output  io_devices_0_ready,
  output  io_devices_0_complete,
  input   io_devices_1_valid,
  output  io_devices_1_ready,
  output  io_devices_1_complete,
  input   io_devices_2_valid,
  output  io_devices_2_ready,
  output  io_devices_2_complete,
  input   io_devices_3_valid,
  output  io_devices_3_ready,
  output  io_devices_3_complete,
  input   io_devices_4_valid,
  output  io_devices_4_ready,
  output  io_devices_4_complete,
  input   io_devices_5_valid,
  output  io_devices_5_ready,
  output  io_devices_5_complete,
  input   io_devices_6_valid,
  output  io_devices_6_ready,
  output  io_devices_6_complete,
  input   io_devices_7_valid,
  output  io_devices_7_ready,
  output  io_devices_7_complete,
  input   io_devices_8_valid,
  output  io_devices_8_ready,
  output  io_devices_8_complete,
  input   io_devices_9_valid,
  output  io_devices_9_ready,
  output  io_devices_9_complete,
  input   io_devices_10_valid,
  output  io_devices_10_ready,
  output  io_devices_10_complete,
  input   io_devices_11_valid,
  output  io_devices_11_ready,
  output  io_devices_11_complete,
  input   io_devices_12_valid,
  output  io_devices_12_ready,
  output  io_devices_12_complete,
  input   io_devices_13_valid,
  output  io_devices_13_ready,
  output  io_devices_13_complete,
  input   io_devices_14_valid,
  output  io_devices_14_ready,
  output  io_devices_14_complete,
  input   io_devices_15_valid,
  output  io_devices_15_ready,
  output  io_devices_15_complete,
  input   io_devices_16_valid,
  output  io_devices_16_ready,
  output  io_devices_16_complete,
  input   io_devices_17_valid,
  output  io_devices_17_ready,
  output  io_devices_17_complete,
  input   io_devices_18_valid,
  output  io_devices_18_ready,
  output  io_devices_18_complete,
  input   io_devices_19_valid,
  output  io_devices_19_ready,
  output  io_devices_19_complete,
  input   io_devices_20_valid,
  output  io_devices_20_ready,
  output  io_devices_20_complete,
  input   io_devices_21_valid,
  output  io_devices_21_ready,
  output  io_devices_21_complete,
  input   io_devices_22_valid,
  output  io_devices_22_ready,
  output  io_devices_22_complete,
  input   io_devices_23_valid,
  output  io_devices_23_ready,
  output  io_devices_23_complete,
  input   io_devices_24_valid,
  output  io_devices_24_ready,
  output  io_devices_24_complete,
  input   io_devices_25_valid,
  output  io_devices_25_ready,
  output  io_devices_25_complete,
  input   io_devices_26_valid,
  output  io_devices_26_ready,
  output  io_devices_26_complete,
  input   io_devices_27_valid,
  output  io_devices_27_ready,
  output  io_devices_27_complete,
  input   io_devices_28_valid,
  output  io_devices_28_ready,
  output  io_devices_28_complete,
  input   io_devices_29_valid,
  output  io_devices_29_ready,
  output  io_devices_29_complete,
  input   io_devices_30_valid,
  output  io_devices_30_ready,
  output  io_devices_30_complete,
  output  io_harts_0,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [11:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data
);
  wire  T_680_0;
  wire  T_680_1;
  wire  T_680_2;
  wire  T_680_3;
  wire  T_680_4;
  wire  T_680_5;
  wire  T_680_6;
  wire  T_680_7;
  wire  T_680_8;
  wire  T_680_9;
  wire  T_680_10;
  wire  T_680_11;
  wire  T_680_12;
  wire  T_680_13;
  wire  T_680_14;
  wire  T_680_15;
  wire  T_680_16;
  wire  T_680_17;
  wire  T_680_18;
  wire  T_680_19;
  wire  T_680_20;
  wire  T_680_21;
  wire  T_680_22;
  wire  T_680_23;
  wire  T_680_24;
  wire  T_680_25;
  wire  T_680_26;
  wire  T_680_27;
  wire  T_680_28;
  wire  T_680_29;
  wire  T_680_30;
  wire  T_680_31;
  wire  priority_0;
  wire  priority_1;
  wire  priority_2;
  wire  priority_3;
  wire  priority_4;
  wire  priority_5;
  wire  priority_6;
  wire  priority_7;
  wire  priority_8;
  wire  priority_9;
  wire  priority_10;
  wire  priority_11;
  wire  priority_12;
  wire  priority_13;
  wire  priority_14;
  wire  priority_15;
  wire  priority_16;
  wire  priority_17;
  wire  priority_18;
  wire  priority_19;
  wire  priority_20;
  wire  priority_21;
  wire  priority_22;
  wire  priority_23;
  wire  priority_24;
  wire  priority_25;
  wire  priority_26;
  wire  priority_27;
  wire  priority_28;
  wire  priority_29;
  wire  priority_30;
  wire  priority_31;
  wire  T_691_0;
  wire  threshold_0;
  wire  T_733_0;
  wire  T_733_1;
  wire  T_733_2;
  wire  T_733_3;
  wire  T_733_4;
  wire  T_733_5;
  wire  T_733_6;
  wire  T_733_7;
  wire  T_733_8;
  wire  T_733_9;
  wire  T_733_10;
  wire  T_733_11;
  wire  T_733_12;
  wire  T_733_13;
  wire  T_733_14;
  wire  T_733_15;
  wire  T_733_16;
  wire  T_733_17;
  wire  T_733_18;
  wire  T_733_19;
  wire  T_733_20;
  wire  T_733_21;
  wire  T_733_22;
  wire  T_733_23;
  wire  T_733_24;
  wire  T_733_25;
  wire  T_733_26;
  wire  T_733_27;
  wire  T_733_28;
  wire  T_733_29;
  wire  T_733_30;
  wire  T_733_31;
  reg  pending_0;
  reg [31:0] GEN_100;
  reg  pending_1;
  reg [31:0] GEN_132;
  reg  pending_2;
  reg [31:0] GEN_133;
  reg  pending_3;
  reg [31:0] GEN_227;
  reg  pending_4;
  reg [31:0] GEN_259;
  reg  pending_5;
  reg [31:0] GEN_260;
  reg  pending_6;
  reg [31:0] GEN_292;
  reg  pending_7;
  reg [31:0] GEN_293;
  reg  pending_8;
  reg [31:0] GEN_325;
  reg  pending_9;
  reg [31:0] GEN_327;
  reg  pending_10;
  reg [31:0] GEN_328;
  reg  pending_11;
  reg [31:0] GEN_360;
  reg  pending_12;
  reg [31:0] GEN_361;
  reg  pending_13;
  reg [31:0] GEN_393;
  reg  pending_14;
  reg [31:0] GEN_394;
  reg  pending_15;
  reg [31:0] GEN_395;
  reg  pending_16;
  reg [31:0] GEN_396;
  reg  pending_17;
  reg [31:0] GEN_397;
  reg  pending_18;
  reg [31:0] GEN_399;
  reg  pending_19;
  reg [31:0] GEN_400;
  reg  pending_20;
  reg [31:0] GEN_402;
  reg  pending_21;
  reg [31:0] GEN_403;
  reg  pending_22;
  reg [31:0] GEN_405;
  reg  pending_23;
  reg [31:0] GEN_406;
  reg  pending_24;
  reg [31:0] GEN_408;
  reg  pending_25;
  reg [31:0] GEN_409;
  reg  pending_26;
  reg [31:0] GEN_411;
  reg  pending_27;
  reg [31:0] GEN_412;
  reg  pending_28;
  reg [31:0] GEN_414;
  reg  pending_29;
  reg [31:0] GEN_415;
  reg  pending_30;
  reg [31:0] GEN_417;
  reg  pending_31;
  reg [31:0] GEN_418;
  reg  enables_0_0;
  reg [31:0] GEN_420;
  reg  enables_0_1;
  reg [31:0] GEN_421;
  reg  enables_0_2;
  reg [31:0] GEN_423;
  reg  enables_0_3;
  reg [31:0] GEN_424;
  reg  enables_0_4;
  reg [31:0] GEN_426;
  reg  enables_0_5;
  reg [31:0] GEN_427;
  reg  enables_0_6;
  reg [31:0] GEN_429;
  reg  enables_0_7;
  reg [31:0] GEN_430;
  reg  enables_0_8;
  reg [31:0] GEN_432;
  reg  enables_0_9;
  reg [31:0] GEN_433;
  reg  enables_0_10;
  reg [31:0] GEN_435;
  reg  enables_0_11;
  reg [31:0] GEN_436;
  reg  enables_0_12;
  reg [31:0] GEN_438;
  reg  enables_0_13;
  reg [31:0] GEN_439;
  reg  enables_0_14;
  reg [31:0] GEN_441;
  reg  enables_0_15;
  reg [31:0] GEN_442;
  reg  enables_0_16;
  reg [31:0] GEN_444;
  reg  enables_0_17;
  reg [31:0] GEN_445;
  reg  enables_0_18;
  reg [31:0] GEN_447;
  reg  enables_0_19;
  reg [31:0] GEN_448;
  reg  enables_0_20;
  reg [31:0] GEN_450;
  reg  enables_0_21;
  reg [31:0] GEN_451;
  reg  enables_0_22;
  reg [31:0] GEN_453;
  reg  enables_0_23;
  reg [31:0] GEN_454;
  reg  enables_0_24;
  reg [31:0] GEN_456;
  reg  enables_0_25;
  reg [31:0] GEN_457;
  reg  enables_0_26;
  reg [31:0] GEN_459;
  reg  enables_0_27;
  reg [31:0] GEN_460;
  reg  enables_0_28;
  reg [31:0] GEN_462;
  reg  enables_0_29;
  reg [31:0] GEN_463;
  reg  enables_0_30;
  reg [31:0] GEN_465;
  reg  enables_0_31;
  reg [31:0] GEN_466;
  wire  T_770;
  wire  GEN_69;
  wire  T_774;
  wire  GEN_70;
  wire  T_778;
  wire  GEN_71;
  wire  T_782;
  wire  GEN_72;
  wire  T_786;
  wire  GEN_73;
  wire  T_790;
  wire  GEN_74;
  wire  T_794;
  wire  GEN_75;
  wire  T_798;
  wire  GEN_76;
  wire  T_802;
  wire  GEN_77;
  wire  T_806;
  wire  GEN_78;
  wire  T_810;
  wire  GEN_79;
  wire  T_814;
  wire  GEN_80;
  wire  T_818;
  wire  GEN_81;
  wire  T_822;
  wire  GEN_82;
  wire  T_826;
  wire  GEN_83;
  wire  T_830;
  wire  GEN_84;
  wire  T_834;
  wire  GEN_85;
  wire  T_838;
  wire  GEN_86;
  wire  T_842;
  wire  GEN_87;
  wire  T_846;
  wire  GEN_88;
  wire  T_850;
  wire  GEN_89;
  wire  T_854;
  wire  GEN_90;
  wire  T_858;
  wire  GEN_91;
  wire  T_862;
  wire  GEN_92;
  wire  T_866;
  wire  GEN_93;
  wire  T_870;
  wire  GEN_94;
  wire  T_874;
  wire  GEN_95;
  wire  T_878;
  wire  GEN_96;
  wire  T_882;
  wire  GEN_97;
  wire  T_886;
  wire  GEN_98;
  wire  T_890;
  wire  GEN_99;
  wire [4:0] maxDevs_0;
  wire  T_900;
  wire [1:0] T_901;
  wire  T_902;
  wire [1:0] T_903;
  wire  T_904;
  wire [1:0] T_905;
  wire  T_906;
  wire [1:0] T_907;
  wire  T_908;
  wire [1:0] T_909;
  wire  T_910;
  wire [1:0] T_911;
  wire  T_912;
  wire [1:0] T_913;
  wire  T_914;
  wire [1:0] T_915;
  wire  T_916;
  wire [1:0] T_917;
  wire  T_918;
  wire [1:0] T_919;
  wire  T_920;
  wire [1:0] T_921;
  wire  T_922;
  wire [1:0] T_923;
  wire  T_924;
  wire [1:0] T_925;
  wire  T_926;
  wire [1:0] T_927;
  wire  T_928;
  wire [1:0] T_929;
  wire  T_930;
  wire [1:0] T_931;
  wire  T_932;
  wire [1:0] T_933;
  wire  T_934;
  wire [1:0] T_935;
  wire  T_936;
  wire [1:0] T_937;
  wire  T_938;
  wire [1:0] T_939;
  wire  T_940;
  wire [1:0] T_941;
  wire  T_942;
  wire [1:0] T_943;
  wire  T_944;
  wire [1:0] T_945;
  wire  T_946;
  wire [1:0] T_947;
  wire  T_948;
  wire [1:0] T_949;
  wire  T_950;
  wire [1:0] T_951;
  wire  T_952;
  wire [1:0] T_953;
  wire  T_954;
  wire [1:0] T_955;
  wire  T_956;
  wire [1:0] T_957;
  wire  T_958;
  wire [1:0] T_959;
  wire  T_960;
  wire [1:0] T_961;
  wire  T_966;
  wire [1:0] T_967;
  wire [1:0] T_969;
  wire  T_970;
  wire  T_971;
  wire  T_974;
  wire [1:0] T_975;
  wire  T_979;
  wire  T_980;
  wire [1:0] T_981;
  wire [1:0] GEN_702;
  wire [2:0] T_983;
  wire [1:0] T_984;
  wire [1:0] T_985;
  wire  T_988;
  wire [1:0] T_989;
  wire  T_993;
  wire  T_996;
  wire [1:0] T_997;
  wire  T_1001;
  wire  T_1002;
  wire [1:0] T_1003;
  wire [1:0] GEN_703;
  wire [2:0] T_1005;
  wire [1:0] T_1006;
  wire [1:0] T_1007;
  wire  T_1008;
  wire [1:0] T_1009;
  wire [2:0] GEN_704;
  wire [3:0] T_1011;
  wire [2:0] T_1012;
  wire [2:0] T_1013;
  wire  T_1016;
  wire [1:0] T_1017;
  wire  T_1021;
  wire  T_1024;
  wire [1:0] T_1025;
  wire  T_1029;
  wire  T_1030;
  wire [1:0] T_1031;
  wire [1:0] GEN_705;
  wire [2:0] T_1033;
  wire [1:0] T_1034;
  wire [1:0] T_1035;
  wire  T_1038;
  wire [1:0] T_1039;
  wire  T_1043;
  wire  T_1046;
  wire [1:0] T_1047;
  wire  T_1051;
  wire  T_1052;
  wire [1:0] T_1053;
  wire [1:0] GEN_706;
  wire [2:0] T_1055;
  wire [1:0] T_1056;
  wire [1:0] T_1057;
  wire  T_1058;
  wire [1:0] T_1059;
  wire [2:0] GEN_707;
  wire [3:0] T_1061;
  wire [2:0] T_1062;
  wire [2:0] T_1063;
  wire  T_1064;
  wire [1:0] T_1065;
  wire [3:0] GEN_708;
  wire [4:0] T_1067;
  wire [3:0] T_1068;
  wire [3:0] T_1069;
  wire  T_1072;
  wire [1:0] T_1073;
  wire  T_1077;
  wire  T_1080;
  wire [1:0] T_1081;
  wire  T_1085;
  wire  T_1086;
  wire [1:0] T_1087;
  wire [1:0] GEN_709;
  wire [2:0] T_1089;
  wire [1:0] T_1090;
  wire [1:0] T_1091;
  wire  T_1094;
  wire [1:0] T_1095;
  wire  T_1099;
  wire  T_1102;
  wire [1:0] T_1103;
  wire  T_1107;
  wire  T_1108;
  wire [1:0] T_1109;
  wire [1:0] GEN_710;
  wire [2:0] T_1111;
  wire [1:0] T_1112;
  wire [1:0] T_1113;
  wire  T_1114;
  wire [1:0] T_1115;
  wire [2:0] GEN_711;
  wire [3:0] T_1117;
  wire [2:0] T_1118;
  wire [2:0] T_1119;
  wire  T_1122;
  wire [1:0] T_1123;
  wire  T_1127;
  wire  T_1130;
  wire [1:0] T_1131;
  wire  T_1135;
  wire  T_1136;
  wire [1:0] T_1137;
  wire [1:0] GEN_712;
  wire [2:0] T_1139;
  wire [1:0] T_1140;
  wire [1:0] T_1141;
  wire  T_1144;
  wire [1:0] T_1145;
  wire  T_1149;
  wire  T_1152;
  wire [1:0] T_1153;
  wire  T_1157;
  wire  T_1158;
  wire [1:0] T_1159;
  wire [1:0] GEN_713;
  wire [2:0] T_1161;
  wire [1:0] T_1162;
  wire [1:0] T_1163;
  wire  T_1164;
  wire [1:0] T_1165;
  wire [2:0] GEN_714;
  wire [3:0] T_1167;
  wire [2:0] T_1168;
  wire [2:0] T_1169;
  wire  T_1170;
  wire [1:0] T_1171;
  wire [3:0] GEN_715;
  wire [4:0] T_1173;
  wire [3:0] T_1174;
  wire [3:0] T_1175;
  wire  T_1176;
  wire [1:0] T_1177;
  wire [4:0] GEN_716;
  wire [5:0] T_1179;
  wire [4:0] T_1180;
  wire [4:0] T_1181;
  reg [4:0] T_1182;
  reg [31:0] GEN_468;
  reg [1:0] T_1183;
  reg [31:0] GEN_469;
  wire [1:0] T_1185;
  wire  T_1186;
  wire  acq_clk;
  wire  acq_reset;
  wire  acq_io_enq_ready;
  wire  acq_io_enq_valid;
  wire [25:0] acq_io_enq_bits_addr_block;
  wire [1:0] acq_io_enq_bits_client_xact_id;
  wire [2:0] acq_io_enq_bits_addr_beat;
  wire  acq_io_enq_bits_is_builtin_type;
  wire [2:0] acq_io_enq_bits_a_type;
  wire [11:0] acq_io_enq_bits_union;
  wire [63:0] acq_io_enq_bits_data;
  wire  acq_io_deq_ready;
  wire  acq_io_deq_valid;
  wire [25:0] acq_io_deq_bits_addr_block;
  wire [1:0] acq_io_deq_bits_client_xact_id;
  wire [2:0] acq_io_deq_bits_addr_beat;
  wire  acq_io_deq_bits_is_builtin_type;
  wire [2:0] acq_io_deq_bits_a_type;
  wire [11:0] acq_io_deq_bits_union;
  wire [63:0] acq_io_deq_bits_data;
  wire  acq_io_count;
  wire  T_1210;
  wire  T_1212;
  wire  T_1213;
  wire  read;
  wire  T_1216;
  wire  T_1217;
  wire  write;
  wire  T_1220;
  wire  T_1221;
  wire  T_1222;
  wire  T_1223;
  wire  T_1225;
  wire [2:0] T_1233_0;
  wire [2:0] T_1233_1;
  wire  T_1235;
  wire  T_1236;
  wire  T_1237;
  wire  T_1238;
  wire [2:0] T_1239;
  wire [2:0] T_1241;
  wire [28:0] T_1242;
  wire [31:0] T_1243;
  wire [25:0] addr;
  wire  hart;
  wire [4:0] GEN_0;
  wire [5:0] T_1245;
  wire [4:0] myMaxDev;
  wire [63:0] rdata;
  wire  T_1251;
  wire  T_1252;
  wire  T_1254;
  wire [1:0] T_1256;
  wire  T_1257;
  wire  T_1258;
  wire [3:0] T_1262;
  wire [3:0] T_1266;
  wire [7:0] T_1267;
  wire  T_1269;
  wire  T_1270;
  wire  T_1274;
  wire [7:0] T_1275;
  wire [7:0] T_1277;
  wire [7:0] T_1278;
  wire  T_1279;
  wire  T_1280;
  wire  T_1281;
  wire  T_1282;
  wire  T_1283;
  wire  T_1284;
  wire  T_1285;
  wire  T_1286;
  wire [7:0] T_1290;
  wire [7:0] T_1294;
  wire [7:0] T_1298;
  wire [7:0] T_1302;
  wire [7:0] T_1306;
  wire [7:0] T_1310;
  wire [7:0] T_1314;
  wire [7:0] T_1318;
  wire [15:0] T_1319;
  wire [15:0] T_1320;
  wire [31:0] T_1321;
  wire [15:0] T_1322;
  wire [15:0] T_1323;
  wire [31:0] T_1324;
  wire [63:0] T_1325;
  wire [63:0] T_1326;
  wire [63:0] T_1403;
  wire [63:0] T_1404;
  wire [63:0] masked_wdata;
  wire  T_1406;
  wire [35:0] T_1409;
  wire  GEN_1;
  wire [36:0] T_1410;
  wire [7:0] T_1412;
  wire [36:0] T_1413;
  wire  T_1414;
  wire  T_1415;
  wire  GEN_2;
  wire  GEN_101;
  wire  GEN_102;
  wire  GEN_103;
  wire  GEN_104;
  wire  GEN_105;
  wire  GEN_106;
  wire  GEN_107;
  wire  GEN_108;
  wire  GEN_109;
  wire  GEN_110;
  wire  GEN_111;
  wire  GEN_112;
  wire  GEN_113;
  wire  GEN_114;
  wire  GEN_115;
  wire  GEN_116;
  wire  GEN_117;
  wire  GEN_118;
  wire  GEN_119;
  wire  GEN_120;
  wire  GEN_121;
  wire  GEN_122;
  wire  GEN_123;
  wire  GEN_124;
  wire  GEN_125;
  wire  GEN_126;
  wire  GEN_127;
  wire  GEN_128;
  wire  GEN_129;
  wire  GEN_130;
  wire  GEN_131;
  wire  GEN_134;
  wire  GEN_135;
  wire  GEN_136;
  wire  GEN_137;
  wire  GEN_138;
  wire  GEN_139;
  wire  GEN_140;
  wire  GEN_141;
  wire  GEN_142;
  wire  GEN_143;
  wire  GEN_144;
  wire  GEN_145;
  wire  GEN_146;
  wire  GEN_147;
  wire  GEN_148;
  wire  GEN_149;
  wire  GEN_150;
  wire  GEN_151;
  wire  GEN_152;
  wire  GEN_153;
  wire  GEN_154;
  wire  GEN_155;
  wire  GEN_156;
  wire  GEN_157;
  wire  GEN_158;
  wire  GEN_159;
  wire  GEN_160;
  wire  GEN_161;
  wire  GEN_162;
  wire  GEN_163;
  wire  GEN_164;
  wire [31:0] T_1447;
  wire [4:0] T_1448;
  wire  GEN_3;
  wire  GEN_717;
  wire  GEN_718;
  wire  GEN_165;
  wire  GEN_720;
  wire  GEN_166;
  wire  GEN_722;
  wire  GEN_167;
  wire  GEN_724;
  wire  GEN_168;
  wire  GEN_726;
  wire  GEN_169;
  wire  GEN_728;
  wire  GEN_170;
  wire  GEN_730;
  wire  GEN_171;
  wire  GEN_732;
  wire  GEN_172;
  wire  GEN_734;
  wire  GEN_173;
  wire  GEN_736;
  wire  GEN_174;
  wire  GEN_738;
  wire  GEN_175;
  wire  GEN_740;
  wire  GEN_176;
  wire  GEN_742;
  wire  GEN_177;
  wire  GEN_744;
  wire  GEN_178;
  wire  GEN_746;
  wire  GEN_179;
  wire  GEN_748;
  wire  GEN_180;
  wire  GEN_750;
  wire  GEN_181;
  wire  GEN_752;
  wire  GEN_182;
  wire  GEN_754;
  wire  GEN_183;
  wire  GEN_756;
  wire  GEN_184;
  wire  GEN_758;
  wire  GEN_185;
  wire  GEN_760;
  wire  GEN_186;
  wire  GEN_762;
  wire  GEN_187;
  wire  GEN_764;
  wire  GEN_188;
  wire  GEN_766;
  wire  GEN_189;
  wire  GEN_768;
  wire  GEN_190;
  wire  GEN_770;
  wire  GEN_191;
  wire  GEN_772;
  wire  GEN_192;
  wire  GEN_774;
  wire  GEN_193;
  wire  GEN_776;
  wire  GEN_194;
  wire  GEN_778;
  wire  GEN_195;
  wire [5:0] T_1450;
  wire [4:0] T_1451;
  wire  GEN_4;
  wire  GEN_196;
  wire  GEN_197;
  wire  GEN_198;
  wire  GEN_199;
  wire  GEN_200;
  wire  GEN_201;
  wire  GEN_202;
  wire  GEN_203;
  wire  GEN_204;
  wire  GEN_205;
  wire  GEN_206;
  wire  GEN_207;
  wire  GEN_208;
  wire  GEN_209;
  wire  GEN_210;
  wire  GEN_211;
  wire  GEN_212;
  wire  GEN_213;
  wire  GEN_214;
  wire  GEN_215;
  wire  GEN_216;
  wire  GEN_217;
  wire  GEN_218;
  wire  GEN_219;
  wire  GEN_220;
  wire  GEN_221;
  wire  GEN_222;
  wire  GEN_223;
  wire  GEN_224;
  wire  GEN_225;
  wire  GEN_226;
  wire  GEN_228;
  wire  GEN_229;
  wire  GEN_230;
  wire  GEN_231;
  wire  GEN_232;
  wire  GEN_233;
  wire  GEN_234;
  wire  GEN_235;
  wire  GEN_236;
  wire  GEN_237;
  wire  GEN_238;
  wire  GEN_239;
  wire  GEN_240;
  wire  GEN_241;
  wire  GEN_242;
  wire  GEN_243;
  wire  GEN_244;
  wire  GEN_245;
  wire  GEN_246;
  wire  GEN_247;
  wire  GEN_248;
  wire  GEN_249;
  wire  GEN_250;
  wire  GEN_251;
  wire  GEN_252;
  wire  GEN_253;
  wire  GEN_254;
  wire  GEN_255;
  wire  GEN_256;
  wire  GEN_257;
  wire  GEN_258;
  wire  GEN_261;
  wire  GEN_262;
  wire  GEN_263;
  wire  GEN_264;
  wire  GEN_265;
  wire  GEN_266;
  wire  GEN_267;
  wire  GEN_268;
  wire  GEN_269;
  wire  GEN_270;
  wire  GEN_271;
  wire  GEN_272;
  wire  GEN_273;
  wire  GEN_274;
  wire  GEN_275;
  wire  GEN_276;
  wire  GEN_277;
  wire  GEN_278;
  wire  GEN_279;
  wire  GEN_280;
  wire  GEN_281;
  wire  GEN_282;
  wire  GEN_283;
  wire  GEN_284;
  wire  GEN_285;
  wire  GEN_286;
  wire  GEN_287;
  wire  GEN_288;
  wire  GEN_289;
  wire  GEN_290;
  wire  GEN_291;
  wire  GEN_294;
  wire  GEN_295;
  wire  GEN_296;
  wire  GEN_297;
  wire  GEN_298;
  wire  GEN_299;
  wire  GEN_300;
  wire  GEN_301;
  wire  GEN_302;
  wire  GEN_303;
  wire  GEN_304;
  wire  GEN_305;
  wire  GEN_306;
  wire  GEN_307;
  wire  GEN_308;
  wire  GEN_309;
  wire  GEN_310;
  wire  GEN_311;
  wire  GEN_312;
  wire  GEN_313;
  wire  GEN_314;
  wire  GEN_315;
  wire  GEN_316;
  wire  GEN_317;
  wire  GEN_318;
  wire  GEN_319;
  wire  GEN_320;
  wire  GEN_321;
  wire  GEN_322;
  wire  GEN_323;
  wire  GEN_324;
  wire [63:0] GEN_326;
  wire  GEN_329;
  wire  GEN_330;
  wire  GEN_331;
  wire  GEN_332;
  wire  GEN_333;
  wire  GEN_334;
  wire  GEN_335;
  wire  GEN_336;
  wire  GEN_337;
  wire  GEN_338;
  wire  GEN_339;
  wire  GEN_340;
  wire  GEN_341;
  wire  GEN_342;
  wire  GEN_343;
  wire  GEN_344;
  wire  GEN_345;
  wire  GEN_346;
  wire  GEN_347;
  wire  GEN_348;
  wire  GEN_349;
  wire  GEN_350;
  wire  GEN_351;
  wire  GEN_352;
  wire  GEN_353;
  wire  GEN_354;
  wire  GEN_355;
  wire  GEN_356;
  wire  GEN_357;
  wire  GEN_358;
  wire  GEN_359;
  wire  GEN_362;
  wire  GEN_363;
  wire  GEN_364;
  wire  GEN_365;
  wire  GEN_366;
  wire  GEN_367;
  wire  GEN_368;
  wire  GEN_369;
  wire  GEN_370;
  wire  GEN_371;
  wire  GEN_372;
  wire  GEN_373;
  wire  GEN_374;
  wire  GEN_375;
  wire  GEN_376;
  wire  GEN_377;
  wire  GEN_378;
  wire  GEN_379;
  wire  GEN_380;
  wire  GEN_381;
  wire  GEN_382;
  wire  GEN_383;
  wire  GEN_384;
  wire  GEN_385;
  wire  GEN_386;
  wire  GEN_387;
  wire  GEN_388;
  wire  GEN_389;
  wire  GEN_390;
  wire  GEN_391;
  wire  GEN_392;
  wire  T_1459;
  wire  T_1461;
  wire  T_1462;
  wire  GEN_5;
  wire  GEN_6;
  wire [1:0] T_1467;
  wire  GEN_7;
  wire  GEN_8;
  wire [1:0] T_1468;
  wire [3:0] T_1469;
  wire  GEN_9;
  wire  GEN_10;
  wire [1:0] T_1470;
  wire  GEN_11;
  wire  GEN_12;
  wire [1:0] T_1471;
  wire [3:0] T_1472;
  wire [7:0] T_1473;
  wire  GEN_13;
  wire  GEN_14;
  wire [1:0] T_1474;
  wire  GEN_15;
  wire  GEN_16;
  wire [1:0] T_1475;
  wire [3:0] T_1476;
  wire  GEN_17;
  wire  GEN_18;
  wire [1:0] T_1477;
  wire  GEN_19;
  wire  GEN_20;
  wire [1:0] T_1478;
  wire [3:0] T_1479;
  wire [7:0] T_1480;
  wire [15:0] T_1481;
  wire  GEN_21;
  wire  GEN_22;
  wire [1:0] T_1482;
  wire  GEN_23;
  wire  GEN_24;
  wire [1:0] T_1483;
  wire [3:0] T_1484;
  wire  GEN_25;
  wire  GEN_26;
  wire [1:0] T_1485;
  wire  GEN_27;
  wire  GEN_28;
  wire [1:0] T_1486;
  wire [3:0] T_1487;
  wire [7:0] T_1488;
  wire  GEN_29;
  wire  GEN_30;
  wire [1:0] T_1489;
  wire  GEN_31;
  wire  GEN_32;
  wire [1:0] T_1490;
  wire [3:0] T_1491;
  wire  GEN_33;
  wire  GEN_34;
  wire [1:0] T_1492;
  wire  GEN_35;
  wire  GEN_36;
  wire [1:0] T_1493;
  wire [3:0] T_1494;
  wire [7:0] T_1495;
  wire [15:0] T_1496;
  wire [31:0] T_1497;
  wire  T_1501;
  wire  GEN_37;
  wire  T_1505;
  wire  GEN_38;
  wire  GEN_398;
  wire  T_1509;
  wire  GEN_39;
  wire  GEN_401;
  wire  T_1513;
  wire  GEN_40;
  wire  GEN_404;
  wire  T_1517;
  wire  GEN_41;
  wire  GEN_407;
  wire  T_1521;
  wire  GEN_42;
  wire  GEN_410;
  wire  T_1525;
  wire  GEN_43;
  wire  GEN_413;
  wire  T_1529;
  wire  GEN_44;
  wire  GEN_416;
  wire  T_1533;
  wire  GEN_45;
  wire  GEN_419;
  wire  T_1537;
  wire  GEN_46;
  wire  GEN_422;
  wire  T_1541;
  wire  GEN_47;
  wire  GEN_425;
  wire  T_1545;
  wire  GEN_48;
  wire  GEN_428;
  wire  T_1549;
  wire  GEN_49;
  wire  GEN_431;
  wire  T_1553;
  wire  GEN_50;
  wire  GEN_434;
  wire  T_1557;
  wire  GEN_51;
  wire  GEN_437;
  wire  T_1561;
  wire  GEN_52;
  wire  GEN_440;
  wire  T_1565;
  wire  GEN_53;
  wire  GEN_443;
  wire  T_1569;
  wire  GEN_54;
  wire  GEN_446;
  wire  T_1573;
  wire  GEN_55;
  wire  GEN_449;
  wire  T_1577;
  wire  GEN_56;
  wire  GEN_452;
  wire  T_1581;
  wire  GEN_57;
  wire  GEN_455;
  wire  T_1585;
  wire  GEN_58;
  wire  GEN_458;
  wire  T_1589;
  wire  GEN_59;
  wire  GEN_461;
  wire  T_1593;
  wire  GEN_60;
  wire  GEN_464;
  wire  T_1597;
  wire  GEN_61;
  wire  GEN_467;
  wire  T_1601;
  wire  GEN_62;
  wire  GEN_470;
  wire  T_1605;
  wire  GEN_63;
  wire  GEN_473;
  wire  T_1609;
  wire  GEN_64;
  wire  GEN_476;
  wire  T_1613;
  wire  GEN_65;
  wire  GEN_479;
  wire  T_1617;
  wire  GEN_66;
  wire  GEN_482;
  wire  T_1621;
  wire  GEN_67;
  wire  GEN_485;
  wire  T_1625;
  wire  GEN_68;
  wire  GEN_488;
  wire [63:0] GEN_521;
  wire [63:0] GEN_619;
  wire  GEN_623;
  wire  GEN_625;
  wire  GEN_627;
  wire  GEN_629;
  wire  GEN_631;
  wire  GEN_633;
  wire  GEN_635;
  wire  GEN_637;
  wire  GEN_639;
  wire  GEN_641;
  wire  GEN_643;
  wire  GEN_645;
  wire  GEN_647;
  wire  GEN_649;
  wire  GEN_651;
  wire  GEN_653;
  wire  GEN_655;
  wire  GEN_657;
  wire  GEN_659;
  wire  GEN_661;
  wire  GEN_663;
  wire  GEN_665;
  wire  GEN_667;
  wire  GEN_669;
  wire  GEN_671;
  wire  GEN_673;
  wire  GEN_675;
  wire  GEN_677;
  wire  GEN_679;
  wire  GEN_681;
  wire  GEN_683;
  wire  T_1627;
  wire  T_1631;
  wire  T_1632;
  wire  T_1633;
  wire [1:0] T_1634;
  wire [1:0] T_1635;
  wire [1:0] T_1636;
  wire [3:0] T_1637;
  wire [1:0] T_1638;
  wire [1:0] T_1639;
  wire [3:0] T_1640;
  wire [7:0] T_1641;
  wire [1:0] T_1642;
  wire [1:0] T_1643;
  wire [3:0] T_1644;
  wire [1:0] T_1645;
  wire [1:0] T_1646;
  wire [3:0] T_1647;
  wire [7:0] T_1648;
  wire [15:0] T_1649;
  wire [1:0] T_1650;
  wire [1:0] T_1651;
  wire [3:0] T_1652;
  wire [1:0] T_1653;
  wire [1:0] T_1654;
  wire [3:0] T_1655;
  wire [7:0] T_1656;
  wire [1:0] T_1657;
  wire [1:0] T_1658;
  wire [3:0] T_1659;
  wire [1:0] T_1660;
  wire [1:0] T_1661;
  wire [3:0] T_1662;
  wire [7:0] T_1663;
  wire [15:0] T_1664;
  wire [31:0] T_1665;
  wire [6:0] GEN_779;
  wire [8:0] T_1667;
  wire [31:0] T_1668;
  wire [63:0] GEN_684;
  wire  T_1675;
  wire  T_1676;
  wire [3:0] T_1677;
  wire  T_1679;
  wire [31:0] T_1681;
  wire [31:0] T_1683;
  wire [63:0] T_1684;
  wire [63:0] GEN_685;
  wire  T_1686;
  wire [31:0] T_1688;
  wire [31:0] T_1690;
  wire [63:0] T_1691;
  wire [63:0] GEN_686;
  wire  T_1693;
  wire [31:0] T_1695;
  wire [31:0] T_1697;
  wire [63:0] T_1698;
  wire [63:0] GEN_687;
  wire  T_1700;
  wire [31:0] T_1702;
  wire [31:0] T_1704;
  wire [63:0] T_1705;
  wire [63:0] GEN_688;
  wire  T_1707;
  wire [31:0] T_1709;
  wire [31:0] T_1711;
  wire [63:0] T_1712;
  wire [63:0] GEN_689;
  wire  T_1714;
  wire [31:0] T_1716;
  wire [31:0] T_1718;
  wire [63:0] T_1719;
  wire [63:0] GEN_690;
  wire  T_1721;
  wire [31:0] T_1723;
  wire [31:0] T_1725;
  wire [63:0] T_1726;
  wire [63:0] GEN_691;
  wire  T_1728;
  wire [31:0] T_1730;
  wire [31:0] T_1732;
  wire [63:0] T_1733;
  wire [63:0] GEN_692;
  wire  T_1735;
  wire [31:0] T_1737;
  wire [31:0] T_1739;
  wire [63:0] T_1740;
  wire [63:0] GEN_693;
  wire  T_1742;
  wire [31:0] T_1744;
  wire [31:0] T_1746;
  wire [63:0] T_1747;
  wire [63:0] GEN_694;
  wire  T_1749;
  wire [31:0] T_1751;
  wire [31:0] T_1753;
  wire [63:0] T_1754;
  wire [63:0] GEN_695;
  wire  T_1756;
  wire [31:0] T_1758;
  wire [31:0] T_1760;
  wire [63:0] T_1761;
  wire [63:0] GEN_696;
  wire  T_1763;
  wire [31:0] T_1765;
  wire [31:0] T_1767;
  wire [63:0] T_1768;
  wire [63:0] GEN_697;
  wire  T_1770;
  wire [31:0] T_1772;
  wire [31:0] T_1774;
  wire [63:0] T_1775;
  wire [63:0] GEN_698;
  wire  T_1777;
  wire [31:0] T_1779;
  wire [31:0] T_1781;
  wire [63:0] T_1782;
  wire [63:0] GEN_699;
  wire  T_1784;
  wire [31:0] T_1786;
  wire [31:0] T_1788;
  wire [63:0] T_1789;
  wire [63:0] GEN_700;
  wire [63:0] GEN_701;
  wire  T_1809;
  wire [2:0] T_1810;
  wire  T_1811;
  wire [2:0] T_1812;
  wire  T_1813;
  wire [2:0] T_1814;
  wire  T_1815;
  wire [2:0] T_1816;
  wire  T_1817;
  wire [2:0] T_1818;
  wire  T_1819;
  wire [2:0] T_1820;
  wire  T_1821;
  wire [2:0] T_1822;
  wire [2:0] T_1847_addr_beat;
  wire [1:0] T_1847_client_xact_id;
  wire  T_1847_manager_xact_id;
  wire  T_1847_is_builtin_type;
  wire [3:0] T_1847_g_type;
  wire [63:0] T_1847_data;
  Queue_8 acq (
    .clk(acq_clk),
    .reset(acq_reset),
    .io_enq_ready(acq_io_enq_ready),
    .io_enq_valid(acq_io_enq_valid),
    .io_enq_bits_addr_block(acq_io_enq_bits_addr_block),
    .io_enq_bits_client_xact_id(acq_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(acq_io_enq_bits_addr_beat),
    .io_enq_bits_is_builtin_type(acq_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(acq_io_enq_bits_a_type),
    .io_enq_bits_union(acq_io_enq_bits_union),
    .io_enq_bits_data(acq_io_enq_bits_data),
    .io_deq_ready(acq_io_deq_ready),
    .io_deq_valid(acq_io_deq_valid),
    .io_deq_bits_addr_block(acq_io_deq_bits_addr_block),
    .io_deq_bits_client_xact_id(acq_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(acq_io_deq_bits_addr_beat),
    .io_deq_bits_is_builtin_type(acq_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(acq_io_deq_bits_a_type),
    .io_deq_bits_union(acq_io_deq_bits_union),
    .io_deq_bits_data(acq_io_deq_bits_data),
    .io_count(acq_io_count)
  );
  assign io_devices_0_ready = T_770;
  assign io_devices_0_complete = GEN_362;
  assign io_devices_1_ready = T_774;
  assign io_devices_1_complete = GEN_363;
  assign io_devices_2_ready = T_778;
  assign io_devices_2_complete = GEN_364;
  assign io_devices_3_ready = T_782;
  assign io_devices_3_complete = GEN_365;
  assign io_devices_4_ready = T_786;
  assign io_devices_4_complete = GEN_366;
  assign io_devices_5_ready = T_790;
  assign io_devices_5_complete = GEN_367;
  assign io_devices_6_ready = T_794;
  assign io_devices_6_complete = GEN_368;
  assign io_devices_7_ready = T_798;
  assign io_devices_7_complete = GEN_369;
  assign io_devices_8_ready = T_802;
  assign io_devices_8_complete = GEN_370;
  assign io_devices_9_ready = T_806;
  assign io_devices_9_complete = GEN_371;
  assign io_devices_10_ready = T_810;
  assign io_devices_10_complete = GEN_372;
  assign io_devices_11_ready = T_814;
  assign io_devices_11_complete = GEN_373;
  assign io_devices_12_ready = T_818;
  assign io_devices_12_complete = GEN_374;
  assign io_devices_13_ready = T_822;
  assign io_devices_13_complete = GEN_375;
  assign io_devices_14_ready = T_826;
  assign io_devices_14_complete = GEN_376;
  assign io_devices_15_ready = T_830;
  assign io_devices_15_complete = GEN_377;
  assign io_devices_16_ready = T_834;
  assign io_devices_16_complete = GEN_378;
  assign io_devices_17_ready = T_838;
  assign io_devices_17_complete = GEN_379;
  assign io_devices_18_ready = T_842;
  assign io_devices_18_complete = GEN_380;
  assign io_devices_19_ready = T_846;
  assign io_devices_19_complete = GEN_381;
  assign io_devices_20_ready = T_850;
  assign io_devices_20_complete = GEN_382;
  assign io_devices_21_ready = T_854;
  assign io_devices_21_complete = GEN_383;
  assign io_devices_22_ready = T_858;
  assign io_devices_22_complete = GEN_384;
  assign io_devices_23_ready = T_862;
  assign io_devices_23_complete = GEN_385;
  assign io_devices_24_ready = T_866;
  assign io_devices_24_complete = GEN_386;
  assign io_devices_25_ready = T_870;
  assign io_devices_25_complete = GEN_387;
  assign io_devices_26_ready = T_874;
  assign io_devices_26_complete = GEN_388;
  assign io_devices_27_ready = T_878;
  assign io_devices_27_complete = GEN_389;
  assign io_devices_28_ready = T_882;
  assign io_devices_28_complete = GEN_390;
  assign io_devices_29_ready = T_886;
  assign io_devices_29_complete = GEN_391;
  assign io_devices_30_ready = T_890;
  assign io_devices_30_complete = GEN_392;
  assign io_harts_0 = T_1186;
  assign io_tl_acquire_ready = acq_io_enq_ready;
  assign io_tl_grant_valid = acq_io_deq_valid;
  assign io_tl_grant_bits_addr_beat = T_1847_addr_beat;
  assign io_tl_grant_bits_client_xact_id = T_1847_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = T_1847_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = T_1847_is_builtin_type;
  assign io_tl_grant_bits_g_type = T_1847_g_type;
  assign io_tl_grant_bits_data = T_1847_data;
  assign T_680_0 = 1'h1;
  assign T_680_1 = 1'h1;
  assign T_680_2 = 1'h1;
  assign T_680_3 = 1'h1;
  assign T_680_4 = 1'h1;
  assign T_680_5 = 1'h1;
  assign T_680_6 = 1'h1;
  assign T_680_7 = 1'h1;
  assign T_680_8 = 1'h1;
  assign T_680_9 = 1'h1;
  assign T_680_10 = 1'h1;
  assign T_680_11 = 1'h1;
  assign T_680_12 = 1'h1;
  assign T_680_13 = 1'h1;
  assign T_680_14 = 1'h1;
  assign T_680_15 = 1'h1;
  assign T_680_16 = 1'h1;
  assign T_680_17 = 1'h1;
  assign T_680_18 = 1'h1;
  assign T_680_19 = 1'h1;
  assign T_680_20 = 1'h1;
  assign T_680_21 = 1'h1;
  assign T_680_22 = 1'h1;
  assign T_680_23 = 1'h1;
  assign T_680_24 = 1'h1;
  assign T_680_25 = 1'h1;
  assign T_680_26 = 1'h1;
  assign T_680_27 = 1'h1;
  assign T_680_28 = 1'h1;
  assign T_680_29 = 1'h1;
  assign T_680_30 = 1'h1;
  assign T_680_31 = 1'h1;
  assign priority_0 = 1'h0;
  assign priority_1 = T_680_1;
  assign priority_2 = T_680_2;
  assign priority_3 = T_680_3;
  assign priority_4 = T_680_4;
  assign priority_5 = T_680_5;
  assign priority_6 = T_680_6;
  assign priority_7 = T_680_7;
  assign priority_8 = T_680_8;
  assign priority_9 = T_680_9;
  assign priority_10 = T_680_10;
  assign priority_11 = T_680_11;
  assign priority_12 = T_680_12;
  assign priority_13 = T_680_13;
  assign priority_14 = T_680_14;
  assign priority_15 = T_680_15;
  assign priority_16 = T_680_16;
  assign priority_17 = T_680_17;
  assign priority_18 = T_680_18;
  assign priority_19 = T_680_19;
  assign priority_20 = T_680_20;
  assign priority_21 = T_680_21;
  assign priority_22 = T_680_22;
  assign priority_23 = T_680_23;
  assign priority_24 = T_680_24;
  assign priority_25 = T_680_25;
  assign priority_26 = T_680_26;
  assign priority_27 = T_680_27;
  assign priority_28 = T_680_28;
  assign priority_29 = T_680_29;
  assign priority_30 = T_680_30;
  assign priority_31 = T_680_31;
  assign T_691_0 = 1'h0;
  assign threshold_0 = T_691_0;
  assign T_733_0 = 1'h0;
  assign T_733_1 = 1'h0;
  assign T_733_2 = 1'h0;
  assign T_733_3 = 1'h0;
  assign T_733_4 = 1'h0;
  assign T_733_5 = 1'h0;
  assign T_733_6 = 1'h0;
  assign T_733_7 = 1'h0;
  assign T_733_8 = 1'h0;
  assign T_733_9 = 1'h0;
  assign T_733_10 = 1'h0;
  assign T_733_11 = 1'h0;
  assign T_733_12 = 1'h0;
  assign T_733_13 = 1'h0;
  assign T_733_14 = 1'h0;
  assign T_733_15 = 1'h0;
  assign T_733_16 = 1'h0;
  assign T_733_17 = 1'h0;
  assign T_733_18 = 1'h0;
  assign T_733_19 = 1'h0;
  assign T_733_20 = 1'h0;
  assign T_733_21 = 1'h0;
  assign T_733_22 = 1'h0;
  assign T_733_23 = 1'h0;
  assign T_733_24 = 1'h0;
  assign T_733_25 = 1'h0;
  assign T_733_26 = 1'h0;
  assign T_733_27 = 1'h0;
  assign T_733_28 = 1'h0;
  assign T_733_29 = 1'h0;
  assign T_733_30 = 1'h0;
  assign T_733_31 = 1'h0;
  assign T_770 = pending_1 == 1'h0;
  assign GEN_69 = io_devices_0_valid ? 1'h1 : pending_1;
  assign T_774 = pending_2 == 1'h0;
  assign GEN_70 = io_devices_1_valid ? 1'h1 : pending_2;
  assign T_778 = pending_3 == 1'h0;
  assign GEN_71 = io_devices_2_valid ? 1'h1 : pending_3;
  assign T_782 = pending_4 == 1'h0;
  assign GEN_72 = io_devices_3_valid ? 1'h1 : pending_4;
  assign T_786 = pending_5 == 1'h0;
  assign GEN_73 = io_devices_4_valid ? 1'h1 : pending_5;
  assign T_790 = pending_6 == 1'h0;
  assign GEN_74 = io_devices_5_valid ? 1'h1 : pending_6;
  assign T_794 = pending_7 == 1'h0;
  assign GEN_75 = io_devices_6_valid ? 1'h1 : pending_7;
  assign T_798 = pending_8 == 1'h0;
  assign GEN_76 = io_devices_7_valid ? 1'h1 : pending_8;
  assign T_802 = pending_9 == 1'h0;
  assign GEN_77 = io_devices_8_valid ? 1'h1 : pending_9;
  assign T_806 = pending_10 == 1'h0;
  assign GEN_78 = io_devices_9_valid ? 1'h1 : pending_10;
  assign T_810 = pending_11 == 1'h0;
  assign GEN_79 = io_devices_10_valid ? 1'h1 : pending_11;
  assign T_814 = pending_12 == 1'h0;
  assign GEN_80 = io_devices_11_valid ? 1'h1 : pending_12;
  assign T_818 = pending_13 == 1'h0;
  assign GEN_81 = io_devices_12_valid ? 1'h1 : pending_13;
  assign T_822 = pending_14 == 1'h0;
  assign GEN_82 = io_devices_13_valid ? 1'h1 : pending_14;
  assign T_826 = pending_15 == 1'h0;
  assign GEN_83 = io_devices_14_valid ? 1'h1 : pending_15;
  assign T_830 = pending_16 == 1'h0;
  assign GEN_84 = io_devices_15_valid ? 1'h1 : pending_16;
  assign T_834 = pending_17 == 1'h0;
  assign GEN_85 = io_devices_16_valid ? 1'h1 : pending_17;
  assign T_838 = pending_18 == 1'h0;
  assign GEN_86 = io_devices_17_valid ? 1'h1 : pending_18;
  assign T_842 = pending_19 == 1'h0;
  assign GEN_87 = io_devices_18_valid ? 1'h1 : pending_19;
  assign T_846 = pending_20 == 1'h0;
  assign GEN_88 = io_devices_19_valid ? 1'h1 : pending_20;
  assign T_850 = pending_21 == 1'h0;
  assign GEN_89 = io_devices_20_valid ? 1'h1 : pending_21;
  assign T_854 = pending_22 == 1'h0;
  assign GEN_90 = io_devices_21_valid ? 1'h1 : pending_22;
  assign T_858 = pending_23 == 1'h0;
  assign GEN_91 = io_devices_22_valid ? 1'h1 : pending_23;
  assign T_862 = pending_24 == 1'h0;
  assign GEN_92 = io_devices_23_valid ? 1'h1 : pending_24;
  assign T_866 = pending_25 == 1'h0;
  assign GEN_93 = io_devices_24_valid ? 1'h1 : pending_25;
  assign T_870 = pending_26 == 1'h0;
  assign GEN_94 = io_devices_25_valid ? 1'h1 : pending_26;
  assign T_874 = pending_27 == 1'h0;
  assign GEN_95 = io_devices_26_valid ? 1'h1 : pending_27;
  assign T_878 = pending_28 == 1'h0;
  assign GEN_96 = io_devices_27_valid ? 1'h1 : pending_28;
  assign T_882 = pending_29 == 1'h0;
  assign GEN_97 = io_devices_28_valid ? 1'h1 : pending_29;
  assign T_886 = pending_30 == 1'h0;
  assign GEN_98 = io_devices_29_valid ? 1'h1 : pending_30;
  assign T_890 = pending_31 == 1'h0;
  assign GEN_99 = io_devices_30_valid ? 1'h1 : pending_31;
  assign maxDevs_0 = T_1182;
  assign T_900 = pending_1 & enables_0_1;
  assign T_901 = {T_900,priority_1};
  assign T_902 = pending_2 & enables_0_2;
  assign T_903 = {T_902,priority_2};
  assign T_904 = pending_3 & enables_0_3;
  assign T_905 = {T_904,priority_3};
  assign T_906 = pending_4 & enables_0_4;
  assign T_907 = {T_906,priority_4};
  assign T_908 = pending_5 & enables_0_5;
  assign T_909 = {T_908,priority_5};
  assign T_910 = pending_6 & enables_0_6;
  assign T_911 = {T_910,priority_6};
  assign T_912 = pending_7 & enables_0_7;
  assign T_913 = {T_912,priority_7};
  assign T_914 = pending_8 & enables_0_8;
  assign T_915 = {T_914,priority_8};
  assign T_916 = pending_9 & enables_0_9;
  assign T_917 = {T_916,priority_9};
  assign T_918 = pending_10 & enables_0_10;
  assign T_919 = {T_918,priority_10};
  assign T_920 = pending_11 & enables_0_11;
  assign T_921 = {T_920,priority_11};
  assign T_922 = pending_12 & enables_0_12;
  assign T_923 = {T_922,priority_12};
  assign T_924 = pending_13 & enables_0_13;
  assign T_925 = {T_924,priority_13};
  assign T_926 = pending_14 & enables_0_14;
  assign T_927 = {T_926,priority_14};
  assign T_928 = pending_15 & enables_0_15;
  assign T_929 = {T_928,priority_15};
  assign T_930 = pending_16 & enables_0_16;
  assign T_931 = {T_930,priority_16};
  assign T_932 = pending_17 & enables_0_17;
  assign T_933 = {T_932,priority_17};
  assign T_934 = pending_18 & enables_0_18;
  assign T_935 = {T_934,priority_18};
  assign T_936 = pending_19 & enables_0_19;
  assign T_937 = {T_936,priority_19};
  assign T_938 = pending_20 & enables_0_20;
  assign T_939 = {T_938,priority_20};
  assign T_940 = pending_21 & enables_0_21;
  assign T_941 = {T_940,priority_21};
  assign T_942 = pending_22 & enables_0_22;
  assign T_943 = {T_942,priority_22};
  assign T_944 = pending_23 & enables_0_23;
  assign T_945 = {T_944,priority_23};
  assign T_946 = pending_24 & enables_0_24;
  assign T_947 = {T_946,priority_24};
  assign T_948 = pending_25 & enables_0_25;
  assign T_949 = {T_948,priority_25};
  assign T_950 = pending_26 & enables_0_26;
  assign T_951 = {T_950,priority_26};
  assign T_952 = pending_27 & enables_0_27;
  assign T_953 = {T_952,priority_27};
  assign T_954 = pending_28 & enables_0_28;
  assign T_955 = {T_954,priority_28};
  assign T_956 = pending_29 & enables_0_29;
  assign T_957 = {T_956,priority_29};
  assign T_958 = pending_30 & enables_0_30;
  assign T_959 = {T_958,priority_30};
  assign T_960 = pending_31 & enables_0_31;
  assign T_961 = {T_960,priority_31};
  assign T_966 = 2'h2 >= T_901;
  assign T_967 = T_966 ? 2'h2 : T_901;
  assign T_969 = 1'h1 + 1'h0;
  assign T_970 = T_969[0:0];
  assign T_971 = T_966 ? 1'h0 : T_970;
  assign T_974 = T_903 >= T_905;
  assign T_975 = T_974 ? T_903 : T_905;
  assign T_979 = T_974 ? 1'h0 : T_970;
  assign T_980 = T_967 >= T_975;
  assign T_981 = T_980 ? T_967 : T_975;
  assign GEN_702 = {{1'd0}, T_979};
  assign T_983 = 2'h2 + GEN_702;
  assign T_984 = T_983[1:0];
  assign T_985 = T_980 ? {{1'd0}, T_971} : T_984;
  assign T_988 = T_907 >= T_909;
  assign T_989 = T_988 ? T_907 : T_909;
  assign T_993 = T_988 ? 1'h0 : T_970;
  assign T_996 = T_911 >= T_913;
  assign T_997 = T_996 ? T_911 : T_913;
  assign T_1001 = T_996 ? 1'h0 : T_970;
  assign T_1002 = T_989 >= T_997;
  assign T_1003 = T_1002 ? T_989 : T_997;
  assign GEN_703 = {{1'd0}, T_1001};
  assign T_1005 = 2'h2 + GEN_703;
  assign T_1006 = T_1005[1:0];
  assign T_1007 = T_1002 ? {{1'd0}, T_993} : T_1006;
  assign T_1008 = T_981 >= T_1003;
  assign T_1009 = T_1008 ? T_981 : T_1003;
  assign GEN_704 = {{1'd0}, T_1007};
  assign T_1011 = 3'h4 + GEN_704;
  assign T_1012 = T_1011[2:0];
  assign T_1013 = T_1008 ? {{1'd0}, T_985} : T_1012;
  assign T_1016 = T_915 >= T_917;
  assign T_1017 = T_1016 ? T_915 : T_917;
  assign T_1021 = T_1016 ? 1'h0 : T_970;
  assign T_1024 = T_919 >= T_921;
  assign T_1025 = T_1024 ? T_919 : T_921;
  assign T_1029 = T_1024 ? 1'h0 : T_970;
  assign T_1030 = T_1017 >= T_1025;
  assign T_1031 = T_1030 ? T_1017 : T_1025;
  assign GEN_705 = {{1'd0}, T_1029};
  assign T_1033 = 2'h2 + GEN_705;
  assign T_1034 = T_1033[1:0];
  assign T_1035 = T_1030 ? {{1'd0}, T_1021} : T_1034;
  assign T_1038 = T_923 >= T_925;
  assign T_1039 = T_1038 ? T_923 : T_925;
  assign T_1043 = T_1038 ? 1'h0 : T_970;
  assign T_1046 = T_927 >= T_929;
  assign T_1047 = T_1046 ? T_927 : T_929;
  assign T_1051 = T_1046 ? 1'h0 : T_970;
  assign T_1052 = T_1039 >= T_1047;
  assign T_1053 = T_1052 ? T_1039 : T_1047;
  assign GEN_706 = {{1'd0}, T_1051};
  assign T_1055 = 2'h2 + GEN_706;
  assign T_1056 = T_1055[1:0];
  assign T_1057 = T_1052 ? {{1'd0}, T_1043} : T_1056;
  assign T_1058 = T_1031 >= T_1053;
  assign T_1059 = T_1058 ? T_1031 : T_1053;
  assign GEN_707 = {{1'd0}, T_1057};
  assign T_1061 = 3'h4 + GEN_707;
  assign T_1062 = T_1061[2:0];
  assign T_1063 = T_1058 ? {{1'd0}, T_1035} : T_1062;
  assign T_1064 = T_1009 >= T_1059;
  assign T_1065 = T_1064 ? T_1009 : T_1059;
  assign GEN_708 = {{1'd0}, T_1063};
  assign T_1067 = 4'h8 + GEN_708;
  assign T_1068 = T_1067[3:0];
  assign T_1069 = T_1064 ? {{1'd0}, T_1013} : T_1068;
  assign T_1072 = T_931 >= T_933;
  assign T_1073 = T_1072 ? T_931 : T_933;
  assign T_1077 = T_1072 ? 1'h0 : T_970;
  assign T_1080 = T_935 >= T_937;
  assign T_1081 = T_1080 ? T_935 : T_937;
  assign T_1085 = T_1080 ? 1'h0 : T_970;
  assign T_1086 = T_1073 >= T_1081;
  assign T_1087 = T_1086 ? T_1073 : T_1081;
  assign GEN_709 = {{1'd0}, T_1085};
  assign T_1089 = 2'h2 + GEN_709;
  assign T_1090 = T_1089[1:0];
  assign T_1091 = T_1086 ? {{1'd0}, T_1077} : T_1090;
  assign T_1094 = T_939 >= T_941;
  assign T_1095 = T_1094 ? T_939 : T_941;
  assign T_1099 = T_1094 ? 1'h0 : T_970;
  assign T_1102 = T_943 >= T_945;
  assign T_1103 = T_1102 ? T_943 : T_945;
  assign T_1107 = T_1102 ? 1'h0 : T_970;
  assign T_1108 = T_1095 >= T_1103;
  assign T_1109 = T_1108 ? T_1095 : T_1103;
  assign GEN_710 = {{1'd0}, T_1107};
  assign T_1111 = 2'h2 + GEN_710;
  assign T_1112 = T_1111[1:0];
  assign T_1113 = T_1108 ? {{1'd0}, T_1099} : T_1112;
  assign T_1114 = T_1087 >= T_1109;
  assign T_1115 = T_1114 ? T_1087 : T_1109;
  assign GEN_711 = {{1'd0}, T_1113};
  assign T_1117 = 3'h4 + GEN_711;
  assign T_1118 = T_1117[2:0];
  assign T_1119 = T_1114 ? {{1'd0}, T_1091} : T_1118;
  assign T_1122 = T_947 >= T_949;
  assign T_1123 = T_1122 ? T_947 : T_949;
  assign T_1127 = T_1122 ? 1'h0 : T_970;
  assign T_1130 = T_951 >= T_953;
  assign T_1131 = T_1130 ? T_951 : T_953;
  assign T_1135 = T_1130 ? 1'h0 : T_970;
  assign T_1136 = T_1123 >= T_1131;
  assign T_1137 = T_1136 ? T_1123 : T_1131;
  assign GEN_712 = {{1'd0}, T_1135};
  assign T_1139 = 2'h2 + GEN_712;
  assign T_1140 = T_1139[1:0];
  assign T_1141 = T_1136 ? {{1'd0}, T_1127} : T_1140;
  assign T_1144 = T_955 >= T_957;
  assign T_1145 = T_1144 ? T_955 : T_957;
  assign T_1149 = T_1144 ? 1'h0 : T_970;
  assign T_1152 = T_959 >= T_961;
  assign T_1153 = T_1152 ? T_959 : T_961;
  assign T_1157 = T_1152 ? 1'h0 : T_970;
  assign T_1158 = T_1145 >= T_1153;
  assign T_1159 = T_1158 ? T_1145 : T_1153;
  assign GEN_713 = {{1'd0}, T_1157};
  assign T_1161 = 2'h2 + GEN_713;
  assign T_1162 = T_1161[1:0];
  assign T_1163 = T_1158 ? {{1'd0}, T_1149} : T_1162;
  assign T_1164 = T_1137 >= T_1159;
  assign T_1165 = T_1164 ? T_1137 : T_1159;
  assign GEN_714 = {{1'd0}, T_1163};
  assign T_1167 = 3'h4 + GEN_714;
  assign T_1168 = T_1167[2:0];
  assign T_1169 = T_1164 ? {{1'd0}, T_1141} : T_1168;
  assign T_1170 = T_1115 >= T_1165;
  assign T_1171 = T_1170 ? T_1115 : T_1165;
  assign GEN_715 = {{1'd0}, T_1169};
  assign T_1173 = 4'h8 + GEN_715;
  assign T_1174 = T_1173[3:0];
  assign T_1175 = T_1170 ? {{1'd0}, T_1119} : T_1174;
  assign T_1176 = T_1065 >= T_1171;
  assign T_1177 = T_1176 ? T_1065 : T_1171;
  assign GEN_716 = {{1'd0}, T_1175};
  assign T_1179 = 5'h10 + GEN_716;
  assign T_1180 = T_1179[4:0];
  assign T_1181 = T_1176 ? {{1'd0}, T_1069} : T_1180;
  assign T_1185 = {1'h1,threshold_0};
  assign T_1186 = T_1183 > T_1185;
  assign acq_clk = clk;
  assign acq_reset = reset;
  assign acq_io_enq_valid = io_tl_acquire_valid;
  assign acq_io_enq_bits_addr_block = io_tl_acquire_bits_addr_block;
  assign acq_io_enq_bits_client_xact_id = io_tl_acquire_bits_client_xact_id;
  assign acq_io_enq_bits_addr_beat = io_tl_acquire_bits_addr_beat;
  assign acq_io_enq_bits_is_builtin_type = io_tl_acquire_bits_is_builtin_type;
  assign acq_io_enq_bits_a_type = io_tl_acquire_bits_a_type;
  assign acq_io_enq_bits_union = io_tl_acquire_bits_union;
  assign acq_io_enq_bits_data = io_tl_acquire_bits_data;
  assign acq_io_deq_ready = io_tl_grant_ready;
  assign T_1210 = acq_io_deq_ready & acq_io_deq_valid;
  assign T_1212 = acq_io_deq_bits_a_type == 3'h0;
  assign T_1213 = acq_io_deq_bits_is_builtin_type & T_1212;
  assign read = T_1210 & T_1213;
  assign T_1216 = acq_io_deq_bits_a_type == 3'h2;
  assign T_1217 = acq_io_deq_bits_is_builtin_type & T_1216;
  assign write = T_1210 & T_1217;
  assign T_1220 = T_1210 == 1'h0;
  assign T_1221 = T_1220 | read;
  assign T_1222 = T_1221 | write;
  assign T_1223 = T_1222 | reset;
  assign T_1225 = T_1223 == 1'h0;
  assign T_1233_0 = 3'h0;
  assign T_1233_1 = 3'h4;
  assign T_1235 = acq_io_deq_bits_a_type == T_1233_0;
  assign T_1236 = acq_io_deq_bits_a_type == T_1233_1;
  assign T_1237 = T_1235 | T_1236;
  assign T_1238 = acq_io_deq_bits_is_builtin_type & T_1237;
  assign T_1239 = acq_io_deq_bits_union[11:9];
  assign T_1241 = T_1238 ? T_1239 : 3'h0;
  assign T_1242 = {acq_io_deq_bits_addr_block,acq_io_deq_bits_addr_beat};
  assign T_1243 = {T_1242,T_1241};
  assign addr = T_1243[25:0];
  assign hart = 1'h0;
  assign GEN_0 = maxDevs_0;
  assign T_1245 = GEN_0 + 5'h0;
  assign myMaxDev = T_1245[4:0];
  assign rdata = GEN_701;
  assign T_1251 = acq_io_deq_bits_a_type == 3'h4;
  assign T_1252 = acq_io_deq_bits_is_builtin_type & T_1251;
  assign T_1254 = T_1239[2];
  assign T_1256 = 2'h1 << T_1254;
  assign T_1257 = T_1256[0];
  assign T_1258 = T_1256[1];
  assign T_1262 = T_1257 ? 4'hf : 4'h0;
  assign T_1266 = T_1258 ? 4'hf : 4'h0;
  assign T_1267 = {T_1266,T_1262};
  assign T_1269 = acq_io_deq_bits_a_type == 3'h3;
  assign T_1270 = acq_io_deq_bits_is_builtin_type & T_1269;
  assign T_1274 = T_1270 | T_1217;
  assign T_1275 = acq_io_deq_bits_union[8:1];
  assign T_1277 = T_1274 ? T_1275 : 8'h0;
  assign T_1278 = T_1252 ? T_1267 : T_1277;
  assign T_1279 = T_1278[0];
  assign T_1280 = T_1278[1];
  assign T_1281 = T_1278[2];
  assign T_1282 = T_1278[3];
  assign T_1283 = T_1278[4];
  assign T_1284 = T_1278[5];
  assign T_1285 = T_1278[6];
  assign T_1286 = T_1278[7];
  assign T_1290 = T_1279 ? 8'hff : 8'h0;
  assign T_1294 = T_1280 ? 8'hff : 8'h0;
  assign T_1298 = T_1281 ? 8'hff : 8'h0;
  assign T_1302 = T_1282 ? 8'hff : 8'h0;
  assign T_1306 = T_1283 ? 8'hff : 8'h0;
  assign T_1310 = T_1284 ? 8'hff : 8'h0;
  assign T_1314 = T_1285 ? 8'hff : 8'h0;
  assign T_1318 = T_1286 ? 8'hff : 8'h0;
  assign T_1319 = {T_1294,T_1290};
  assign T_1320 = {T_1302,T_1298};
  assign T_1321 = {T_1320,T_1319};
  assign T_1322 = {T_1310,T_1306};
  assign T_1323 = {T_1318,T_1314};
  assign T_1324 = {T_1323,T_1322};
  assign T_1325 = {T_1324,T_1321};
  assign T_1326 = acq_io_deq_bits_data & T_1325;
  assign T_1403 = ~ T_1325;
  assign T_1404 = rdata & T_1403;
  assign masked_wdata = T_1326 | T_1404;
  assign T_1406 = addr >= 26'h200000;
  assign T_1409 = {myMaxDev,31'h0};
  assign GEN_1 = threshold_0;
  assign T_1410 = {T_1409,GEN_1};
  assign T_1412 = 7'h0 * 7'h40;
  assign T_1413 = T_1410 >> T_1412;
  assign T_1414 = addr[2];
  assign T_1415 = read & T_1414;
  assign GEN_2 = 1'h0;
  assign GEN_101 = 5'h1 == myMaxDev ? GEN_2 : GEN_69;
  assign GEN_102 = 5'h2 == myMaxDev ? GEN_2 : GEN_70;
  assign GEN_103 = 5'h3 == myMaxDev ? GEN_2 : GEN_71;
  assign GEN_104 = 5'h4 == myMaxDev ? GEN_2 : GEN_72;
  assign GEN_105 = 5'h5 == myMaxDev ? GEN_2 : GEN_73;
  assign GEN_106 = 5'h6 == myMaxDev ? GEN_2 : GEN_74;
  assign GEN_107 = 5'h7 == myMaxDev ? GEN_2 : GEN_75;
  assign GEN_108 = 5'h8 == myMaxDev ? GEN_2 : GEN_76;
  assign GEN_109 = 5'h9 == myMaxDev ? GEN_2 : GEN_77;
  assign GEN_110 = 5'ha == myMaxDev ? GEN_2 : GEN_78;
  assign GEN_111 = 5'hb == myMaxDev ? GEN_2 : GEN_79;
  assign GEN_112 = 5'hc == myMaxDev ? GEN_2 : GEN_80;
  assign GEN_113 = 5'hd == myMaxDev ? GEN_2 : GEN_81;
  assign GEN_114 = 5'he == myMaxDev ? GEN_2 : GEN_82;
  assign GEN_115 = 5'hf == myMaxDev ? GEN_2 : GEN_83;
  assign GEN_116 = 5'h10 == myMaxDev ? GEN_2 : GEN_84;
  assign GEN_117 = 5'h11 == myMaxDev ? GEN_2 : GEN_85;
  assign GEN_118 = 5'h12 == myMaxDev ? GEN_2 : GEN_86;
  assign GEN_119 = 5'h13 == myMaxDev ? GEN_2 : GEN_87;
  assign GEN_120 = 5'h14 == myMaxDev ? GEN_2 : GEN_88;
  assign GEN_121 = 5'h15 == myMaxDev ? GEN_2 : GEN_89;
  assign GEN_122 = 5'h16 == myMaxDev ? GEN_2 : GEN_90;
  assign GEN_123 = 5'h17 == myMaxDev ? GEN_2 : GEN_91;
  assign GEN_124 = 5'h18 == myMaxDev ? GEN_2 : GEN_92;
  assign GEN_125 = 5'h19 == myMaxDev ? GEN_2 : GEN_93;
  assign GEN_126 = 5'h1a == myMaxDev ? GEN_2 : GEN_94;
  assign GEN_127 = 5'h1b == myMaxDev ? GEN_2 : GEN_95;
  assign GEN_128 = 5'h1c == myMaxDev ? GEN_2 : GEN_96;
  assign GEN_129 = 5'h1d == myMaxDev ? GEN_2 : GEN_97;
  assign GEN_130 = 5'h1e == myMaxDev ? GEN_2 : GEN_98;
  assign GEN_131 = 5'h1f == myMaxDev ? GEN_2 : GEN_99;
  assign GEN_134 = T_1415 ? GEN_101 : GEN_69;
  assign GEN_135 = T_1415 ? GEN_102 : GEN_70;
  assign GEN_136 = T_1415 ? GEN_103 : GEN_71;
  assign GEN_137 = T_1415 ? GEN_104 : GEN_72;
  assign GEN_138 = T_1415 ? GEN_105 : GEN_73;
  assign GEN_139 = T_1415 ? GEN_106 : GEN_74;
  assign GEN_140 = T_1415 ? GEN_107 : GEN_75;
  assign GEN_141 = T_1415 ? GEN_108 : GEN_76;
  assign GEN_142 = T_1415 ? GEN_109 : GEN_77;
  assign GEN_143 = T_1415 ? GEN_110 : GEN_78;
  assign GEN_144 = T_1415 ? GEN_111 : GEN_79;
  assign GEN_145 = T_1415 ? GEN_112 : GEN_80;
  assign GEN_146 = T_1415 ? GEN_113 : GEN_81;
  assign GEN_147 = T_1415 ? GEN_114 : GEN_82;
  assign GEN_148 = T_1415 ? GEN_115 : GEN_83;
  assign GEN_149 = T_1415 ? GEN_116 : GEN_84;
  assign GEN_150 = T_1415 ? GEN_117 : GEN_85;
  assign GEN_151 = T_1415 ? GEN_118 : GEN_86;
  assign GEN_152 = T_1415 ? GEN_119 : GEN_87;
  assign GEN_153 = T_1415 ? GEN_120 : GEN_88;
  assign GEN_154 = T_1415 ? GEN_121 : GEN_89;
  assign GEN_155 = T_1415 ? GEN_122 : GEN_90;
  assign GEN_156 = T_1415 ? GEN_123 : GEN_91;
  assign GEN_157 = T_1415 ? GEN_124 : GEN_92;
  assign GEN_158 = T_1415 ? GEN_125 : GEN_93;
  assign GEN_159 = T_1415 ? GEN_126 : GEN_94;
  assign GEN_160 = T_1415 ? GEN_127 : GEN_95;
  assign GEN_161 = T_1415 ? GEN_128 : GEN_96;
  assign GEN_162 = T_1415 ? GEN_129 : GEN_97;
  assign GEN_163 = T_1415 ? GEN_130 : GEN_98;
  assign GEN_164 = T_1415 ? GEN_131 : GEN_99;
  assign T_1447 = acq_io_deq_bits_data[63:32];
  assign T_1448 = T_1447[4:0];
  assign GEN_3 = GEN_195;
  assign GEN_717 = 1'h0 == hart;
  assign GEN_718 = 5'h1 == T_1448;
  assign GEN_165 = GEN_717 & GEN_718 ? enables_0_1 : enables_0_0;
  assign GEN_720 = 5'h2 == T_1448;
  assign GEN_166 = GEN_717 & GEN_720 ? enables_0_2 : GEN_165;
  assign GEN_722 = 5'h3 == T_1448;
  assign GEN_167 = GEN_717 & GEN_722 ? enables_0_3 : GEN_166;
  assign GEN_724 = 5'h4 == T_1448;
  assign GEN_168 = GEN_717 & GEN_724 ? enables_0_4 : GEN_167;
  assign GEN_726 = 5'h5 == T_1448;
  assign GEN_169 = GEN_717 & GEN_726 ? enables_0_5 : GEN_168;
  assign GEN_728 = 5'h6 == T_1448;
  assign GEN_170 = GEN_717 & GEN_728 ? enables_0_6 : GEN_169;
  assign GEN_730 = 5'h7 == T_1448;
  assign GEN_171 = GEN_717 & GEN_730 ? enables_0_7 : GEN_170;
  assign GEN_732 = 5'h8 == T_1448;
  assign GEN_172 = GEN_717 & GEN_732 ? enables_0_8 : GEN_171;
  assign GEN_734 = 5'h9 == T_1448;
  assign GEN_173 = GEN_717 & GEN_734 ? enables_0_9 : GEN_172;
  assign GEN_736 = 5'ha == T_1448;
  assign GEN_174 = GEN_717 & GEN_736 ? enables_0_10 : GEN_173;
  assign GEN_738 = 5'hb == T_1448;
  assign GEN_175 = GEN_717 & GEN_738 ? enables_0_11 : GEN_174;
  assign GEN_740 = 5'hc == T_1448;
  assign GEN_176 = GEN_717 & GEN_740 ? enables_0_12 : GEN_175;
  assign GEN_742 = 5'hd == T_1448;
  assign GEN_177 = GEN_717 & GEN_742 ? enables_0_13 : GEN_176;
  assign GEN_744 = 5'he == T_1448;
  assign GEN_178 = GEN_717 & GEN_744 ? enables_0_14 : GEN_177;
  assign GEN_746 = 5'hf == T_1448;
  assign GEN_179 = GEN_717 & GEN_746 ? enables_0_15 : GEN_178;
  assign GEN_748 = 5'h10 == T_1448;
  assign GEN_180 = GEN_717 & GEN_748 ? enables_0_16 : GEN_179;
  assign GEN_750 = 5'h11 == T_1448;
  assign GEN_181 = GEN_717 & GEN_750 ? enables_0_17 : GEN_180;
  assign GEN_752 = 5'h12 == T_1448;
  assign GEN_182 = GEN_717 & GEN_752 ? enables_0_18 : GEN_181;
  assign GEN_754 = 5'h13 == T_1448;
  assign GEN_183 = GEN_717 & GEN_754 ? enables_0_19 : GEN_182;
  assign GEN_756 = 5'h14 == T_1448;
  assign GEN_184 = GEN_717 & GEN_756 ? enables_0_20 : GEN_183;
  assign GEN_758 = 5'h15 == T_1448;
  assign GEN_185 = GEN_717 & GEN_758 ? enables_0_21 : GEN_184;
  assign GEN_760 = 5'h16 == T_1448;
  assign GEN_186 = GEN_717 & GEN_760 ? enables_0_22 : GEN_185;
  assign GEN_762 = 5'h17 == T_1448;
  assign GEN_187 = GEN_717 & GEN_762 ? enables_0_23 : GEN_186;
  assign GEN_764 = 5'h18 == T_1448;
  assign GEN_188 = GEN_717 & GEN_764 ? enables_0_24 : GEN_187;
  assign GEN_766 = 5'h19 == T_1448;
  assign GEN_189 = GEN_717 & GEN_766 ? enables_0_25 : GEN_188;
  assign GEN_768 = 5'h1a == T_1448;
  assign GEN_190 = GEN_717 & GEN_768 ? enables_0_26 : GEN_189;
  assign GEN_770 = 5'h1b == T_1448;
  assign GEN_191 = GEN_717 & GEN_770 ? enables_0_27 : GEN_190;
  assign GEN_772 = 5'h1c == T_1448;
  assign GEN_192 = GEN_717 & GEN_772 ? enables_0_28 : GEN_191;
  assign GEN_774 = 5'h1d == T_1448;
  assign GEN_193 = GEN_717 & GEN_774 ? enables_0_29 : GEN_192;
  assign GEN_776 = 5'h1e == T_1448;
  assign GEN_194 = GEN_717 & GEN_776 ? enables_0_30 : GEN_193;
  assign GEN_778 = 5'h1f == T_1448;
  assign GEN_195 = GEN_717 & GEN_778 ? enables_0_31 : GEN_194;
  assign T_1450 = T_1448 - 5'h1;
  assign T_1451 = T_1450[4:0];
  assign GEN_4 = 1'h1;
  assign GEN_196 = 5'h0 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_197 = 5'h1 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_198 = 5'h2 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_199 = 5'h3 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_200 = 5'h4 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_201 = 5'h5 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_202 = 5'h6 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_203 = 5'h7 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_204 = 5'h8 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_205 = 5'h9 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_206 = 5'ha == T_1451 ? GEN_4 : 1'h0;
  assign GEN_207 = 5'hb == T_1451 ? GEN_4 : 1'h0;
  assign GEN_208 = 5'hc == T_1451 ? GEN_4 : 1'h0;
  assign GEN_209 = 5'hd == T_1451 ? GEN_4 : 1'h0;
  assign GEN_210 = 5'he == T_1451 ? GEN_4 : 1'h0;
  assign GEN_211 = 5'hf == T_1451 ? GEN_4 : 1'h0;
  assign GEN_212 = 5'h10 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_213 = 5'h11 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_214 = 5'h12 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_215 = 5'h13 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_216 = 5'h14 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_217 = 5'h15 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_218 = 5'h16 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_219 = 5'h17 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_220 = 5'h18 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_221 = 5'h19 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_222 = 5'h1a == T_1451 ? GEN_4 : 1'h0;
  assign GEN_223 = 5'h1b == T_1451 ? GEN_4 : 1'h0;
  assign GEN_224 = 5'h1c == T_1451 ? GEN_4 : 1'h0;
  assign GEN_225 = 5'h1d == T_1451 ? GEN_4 : 1'h0;
  assign GEN_226 = 5'h1e == T_1451 ? GEN_4 : 1'h0;
  assign GEN_228 = GEN_3 ? GEN_196 : 1'h0;
  assign GEN_229 = GEN_3 ? GEN_197 : 1'h0;
  assign GEN_230 = GEN_3 ? GEN_198 : 1'h0;
  assign GEN_231 = GEN_3 ? GEN_199 : 1'h0;
  assign GEN_232 = GEN_3 ? GEN_200 : 1'h0;
  assign GEN_233 = GEN_3 ? GEN_201 : 1'h0;
  assign GEN_234 = GEN_3 ? GEN_202 : 1'h0;
  assign GEN_235 = GEN_3 ? GEN_203 : 1'h0;
  assign GEN_236 = GEN_3 ? GEN_204 : 1'h0;
  assign GEN_237 = GEN_3 ? GEN_205 : 1'h0;
  assign GEN_238 = GEN_3 ? GEN_206 : 1'h0;
  assign GEN_239 = GEN_3 ? GEN_207 : 1'h0;
  assign GEN_240 = GEN_3 ? GEN_208 : 1'h0;
  assign GEN_241 = GEN_3 ? GEN_209 : 1'h0;
  assign GEN_242 = GEN_3 ? GEN_210 : 1'h0;
  assign GEN_243 = GEN_3 ? GEN_211 : 1'h0;
  assign GEN_244 = GEN_3 ? GEN_212 : 1'h0;
  assign GEN_245 = GEN_3 ? GEN_213 : 1'h0;
  assign GEN_246 = GEN_3 ? GEN_214 : 1'h0;
  assign GEN_247 = GEN_3 ? GEN_215 : 1'h0;
  assign GEN_248 = GEN_3 ? GEN_216 : 1'h0;
  assign GEN_249 = GEN_3 ? GEN_217 : 1'h0;
  assign GEN_250 = GEN_3 ? GEN_218 : 1'h0;
  assign GEN_251 = GEN_3 ? GEN_219 : 1'h0;
  assign GEN_252 = GEN_3 ? GEN_220 : 1'h0;
  assign GEN_253 = GEN_3 ? GEN_221 : 1'h0;
  assign GEN_254 = GEN_3 ? GEN_222 : 1'h0;
  assign GEN_255 = GEN_3 ? GEN_223 : 1'h0;
  assign GEN_256 = GEN_3 ? GEN_224 : 1'h0;
  assign GEN_257 = GEN_3 ? GEN_225 : 1'h0;
  assign GEN_258 = GEN_3 ? GEN_226 : 1'h0;
  assign GEN_261 = T_1283 ? GEN_228 : 1'h0;
  assign GEN_262 = T_1283 ? GEN_229 : 1'h0;
  assign GEN_263 = T_1283 ? GEN_230 : 1'h0;
  assign GEN_264 = T_1283 ? GEN_231 : 1'h0;
  assign GEN_265 = T_1283 ? GEN_232 : 1'h0;
  assign GEN_266 = T_1283 ? GEN_233 : 1'h0;
  assign GEN_267 = T_1283 ? GEN_234 : 1'h0;
  assign GEN_268 = T_1283 ? GEN_235 : 1'h0;
  assign GEN_269 = T_1283 ? GEN_236 : 1'h0;
  assign GEN_270 = T_1283 ? GEN_237 : 1'h0;
  assign GEN_271 = T_1283 ? GEN_238 : 1'h0;
  assign GEN_272 = T_1283 ? GEN_239 : 1'h0;
  assign GEN_273 = T_1283 ? GEN_240 : 1'h0;
  assign GEN_274 = T_1283 ? GEN_241 : 1'h0;
  assign GEN_275 = T_1283 ? GEN_242 : 1'h0;
  assign GEN_276 = T_1283 ? GEN_243 : 1'h0;
  assign GEN_277 = T_1283 ? GEN_244 : 1'h0;
  assign GEN_278 = T_1283 ? GEN_245 : 1'h0;
  assign GEN_279 = T_1283 ? GEN_246 : 1'h0;
  assign GEN_280 = T_1283 ? GEN_247 : 1'h0;
  assign GEN_281 = T_1283 ? GEN_248 : 1'h0;
  assign GEN_282 = T_1283 ? GEN_249 : 1'h0;
  assign GEN_283 = T_1283 ? GEN_250 : 1'h0;
  assign GEN_284 = T_1283 ? GEN_251 : 1'h0;
  assign GEN_285 = T_1283 ? GEN_252 : 1'h0;
  assign GEN_286 = T_1283 ? GEN_253 : 1'h0;
  assign GEN_287 = T_1283 ? GEN_254 : 1'h0;
  assign GEN_288 = T_1283 ? GEN_255 : 1'h0;
  assign GEN_289 = T_1283 ? GEN_256 : 1'h0;
  assign GEN_290 = T_1283 ? GEN_257 : 1'h0;
  assign GEN_291 = T_1283 ? GEN_258 : 1'h0;
  assign GEN_294 = write ? GEN_261 : 1'h0;
  assign GEN_295 = write ? GEN_262 : 1'h0;
  assign GEN_296 = write ? GEN_263 : 1'h0;
  assign GEN_297 = write ? GEN_264 : 1'h0;
  assign GEN_298 = write ? GEN_265 : 1'h0;
  assign GEN_299 = write ? GEN_266 : 1'h0;
  assign GEN_300 = write ? GEN_267 : 1'h0;
  assign GEN_301 = write ? GEN_268 : 1'h0;
  assign GEN_302 = write ? GEN_269 : 1'h0;
  assign GEN_303 = write ? GEN_270 : 1'h0;
  assign GEN_304 = write ? GEN_271 : 1'h0;
  assign GEN_305 = write ? GEN_272 : 1'h0;
  assign GEN_306 = write ? GEN_273 : 1'h0;
  assign GEN_307 = write ? GEN_274 : 1'h0;
  assign GEN_308 = write ? GEN_275 : 1'h0;
  assign GEN_309 = write ? GEN_276 : 1'h0;
  assign GEN_310 = write ? GEN_277 : 1'h0;
  assign GEN_311 = write ? GEN_278 : 1'h0;
  assign GEN_312 = write ? GEN_279 : 1'h0;
  assign GEN_313 = write ? GEN_280 : 1'h0;
  assign GEN_314 = write ? GEN_281 : 1'h0;
  assign GEN_315 = write ? GEN_282 : 1'h0;
  assign GEN_316 = write ? GEN_283 : 1'h0;
  assign GEN_317 = write ? GEN_284 : 1'h0;
  assign GEN_318 = write ? GEN_285 : 1'h0;
  assign GEN_319 = write ? GEN_286 : 1'h0;
  assign GEN_320 = write ? GEN_287 : 1'h0;
  assign GEN_321 = write ? GEN_288 : 1'h0;
  assign GEN_322 = write ? GEN_289 : 1'h0;
  assign GEN_323 = write ? GEN_290 : 1'h0;
  assign GEN_324 = write ? GEN_291 : 1'h0;
  assign GEN_326 = T_1406 ? {{27'd0}, T_1413} : 64'h0;
  assign GEN_329 = T_1406 ? GEN_134 : GEN_69;
  assign GEN_330 = T_1406 ? GEN_135 : GEN_70;
  assign GEN_331 = T_1406 ? GEN_136 : GEN_71;
  assign GEN_332 = T_1406 ? GEN_137 : GEN_72;
  assign GEN_333 = T_1406 ? GEN_138 : GEN_73;
  assign GEN_334 = T_1406 ? GEN_139 : GEN_74;
  assign GEN_335 = T_1406 ? GEN_140 : GEN_75;
  assign GEN_336 = T_1406 ? GEN_141 : GEN_76;
  assign GEN_337 = T_1406 ? GEN_142 : GEN_77;
  assign GEN_338 = T_1406 ? GEN_143 : GEN_78;
  assign GEN_339 = T_1406 ? GEN_144 : GEN_79;
  assign GEN_340 = T_1406 ? GEN_145 : GEN_80;
  assign GEN_341 = T_1406 ? GEN_146 : GEN_81;
  assign GEN_342 = T_1406 ? GEN_147 : GEN_82;
  assign GEN_343 = T_1406 ? GEN_148 : GEN_83;
  assign GEN_344 = T_1406 ? GEN_149 : GEN_84;
  assign GEN_345 = T_1406 ? GEN_150 : GEN_85;
  assign GEN_346 = T_1406 ? GEN_151 : GEN_86;
  assign GEN_347 = T_1406 ? GEN_152 : GEN_87;
  assign GEN_348 = T_1406 ? GEN_153 : GEN_88;
  assign GEN_349 = T_1406 ? GEN_154 : GEN_89;
  assign GEN_350 = T_1406 ? GEN_155 : GEN_90;
  assign GEN_351 = T_1406 ? GEN_156 : GEN_91;
  assign GEN_352 = T_1406 ? GEN_157 : GEN_92;
  assign GEN_353 = T_1406 ? GEN_158 : GEN_93;
  assign GEN_354 = T_1406 ? GEN_159 : GEN_94;
  assign GEN_355 = T_1406 ? GEN_160 : GEN_95;
  assign GEN_356 = T_1406 ? GEN_161 : GEN_96;
  assign GEN_357 = T_1406 ? GEN_162 : GEN_97;
  assign GEN_358 = T_1406 ? GEN_163 : GEN_98;
  assign GEN_359 = T_1406 ? GEN_164 : GEN_99;
  assign GEN_362 = T_1406 ? GEN_294 : 1'h0;
  assign GEN_363 = T_1406 ? GEN_295 : 1'h0;
  assign GEN_364 = T_1406 ? GEN_296 : 1'h0;
  assign GEN_365 = T_1406 ? GEN_297 : 1'h0;
  assign GEN_366 = T_1406 ? GEN_298 : 1'h0;
  assign GEN_367 = T_1406 ? GEN_299 : 1'h0;
  assign GEN_368 = T_1406 ? GEN_300 : 1'h0;
  assign GEN_369 = T_1406 ? GEN_301 : 1'h0;
  assign GEN_370 = T_1406 ? GEN_302 : 1'h0;
  assign GEN_371 = T_1406 ? GEN_303 : 1'h0;
  assign GEN_372 = T_1406 ? GEN_304 : 1'h0;
  assign GEN_373 = T_1406 ? GEN_305 : 1'h0;
  assign GEN_374 = T_1406 ? GEN_306 : 1'h0;
  assign GEN_375 = T_1406 ? GEN_307 : 1'h0;
  assign GEN_376 = T_1406 ? GEN_308 : 1'h0;
  assign GEN_377 = T_1406 ? GEN_309 : 1'h0;
  assign GEN_378 = T_1406 ? GEN_310 : 1'h0;
  assign GEN_379 = T_1406 ? GEN_311 : 1'h0;
  assign GEN_380 = T_1406 ? GEN_312 : 1'h0;
  assign GEN_381 = T_1406 ? GEN_313 : 1'h0;
  assign GEN_382 = T_1406 ? GEN_314 : 1'h0;
  assign GEN_383 = T_1406 ? GEN_315 : 1'h0;
  assign GEN_384 = T_1406 ? GEN_316 : 1'h0;
  assign GEN_385 = T_1406 ? GEN_317 : 1'h0;
  assign GEN_386 = T_1406 ? GEN_318 : 1'h0;
  assign GEN_387 = T_1406 ? GEN_319 : 1'h0;
  assign GEN_388 = T_1406 ? GEN_320 : 1'h0;
  assign GEN_389 = T_1406 ? GEN_321 : 1'h0;
  assign GEN_390 = T_1406 ? GEN_322 : 1'h0;
  assign GEN_391 = T_1406 ? GEN_323 : 1'h0;
  assign GEN_392 = T_1406 ? GEN_324 : 1'h0;
  assign T_1459 = addr >= 26'h2000;
  assign T_1461 = T_1406 == 1'h0;
  assign T_1462 = T_1461 & T_1459;
  assign GEN_5 = enables_0_1;
  assign GEN_6 = enables_0_0;
  assign T_1467 = {GEN_5,GEN_6};
  assign GEN_7 = enables_0_3;
  assign GEN_8 = enables_0_2;
  assign T_1468 = {GEN_7,GEN_8};
  assign T_1469 = {T_1468,T_1467};
  assign GEN_9 = enables_0_5;
  assign GEN_10 = enables_0_4;
  assign T_1470 = {GEN_9,GEN_10};
  assign GEN_11 = enables_0_7;
  assign GEN_12 = enables_0_6;
  assign T_1471 = {GEN_11,GEN_12};
  assign T_1472 = {T_1471,T_1470};
  assign T_1473 = {T_1472,T_1469};
  assign GEN_13 = enables_0_9;
  assign GEN_14 = enables_0_8;
  assign T_1474 = {GEN_13,GEN_14};
  assign GEN_15 = enables_0_11;
  assign GEN_16 = enables_0_10;
  assign T_1475 = {GEN_15,GEN_16};
  assign T_1476 = {T_1475,T_1474};
  assign GEN_17 = enables_0_13;
  assign GEN_18 = enables_0_12;
  assign T_1477 = {GEN_17,GEN_18};
  assign GEN_19 = enables_0_15;
  assign GEN_20 = enables_0_14;
  assign T_1478 = {GEN_19,GEN_20};
  assign T_1479 = {T_1478,T_1477};
  assign T_1480 = {T_1479,T_1476};
  assign T_1481 = {T_1480,T_1473};
  assign GEN_21 = enables_0_17;
  assign GEN_22 = enables_0_16;
  assign T_1482 = {GEN_21,GEN_22};
  assign GEN_23 = enables_0_19;
  assign GEN_24 = enables_0_18;
  assign T_1483 = {GEN_23,GEN_24};
  assign T_1484 = {T_1483,T_1482};
  assign GEN_25 = enables_0_21;
  assign GEN_26 = enables_0_20;
  assign T_1485 = {GEN_25,GEN_26};
  assign GEN_27 = enables_0_23;
  assign GEN_28 = enables_0_22;
  assign T_1486 = {GEN_27,GEN_28};
  assign T_1487 = {T_1486,T_1485};
  assign T_1488 = {T_1487,T_1484};
  assign GEN_29 = enables_0_25;
  assign GEN_30 = enables_0_24;
  assign T_1489 = {GEN_29,GEN_30};
  assign GEN_31 = enables_0_27;
  assign GEN_32 = enables_0_26;
  assign T_1490 = {GEN_31,GEN_32};
  assign T_1491 = {T_1490,T_1489};
  assign GEN_33 = enables_0_29;
  assign GEN_34 = enables_0_28;
  assign T_1492 = {GEN_33,GEN_34};
  assign GEN_35 = enables_0_31;
  assign GEN_36 = enables_0_30;
  assign T_1493 = {GEN_35,GEN_36};
  assign T_1494 = {T_1493,T_1492};
  assign T_1495 = {T_1494,T_1491};
  assign T_1496 = {T_1495,T_1488};
  assign T_1497 = {T_1496,T_1481};
  assign T_1501 = masked_wdata[0];
  assign GEN_37 = T_1501;
  assign T_1505 = masked_wdata[1];
  assign GEN_38 = T_1505;
  assign GEN_398 = write ? GEN_38 : enables_0_1;
  assign T_1509 = masked_wdata[2];
  assign GEN_39 = T_1509;
  assign GEN_401 = write ? GEN_39 : enables_0_2;
  assign T_1513 = masked_wdata[3];
  assign GEN_40 = T_1513;
  assign GEN_404 = write ? GEN_40 : enables_0_3;
  assign T_1517 = masked_wdata[4];
  assign GEN_41 = T_1517;
  assign GEN_407 = write ? GEN_41 : enables_0_4;
  assign T_1521 = masked_wdata[5];
  assign GEN_42 = T_1521;
  assign GEN_410 = write ? GEN_42 : enables_0_5;
  assign T_1525 = masked_wdata[6];
  assign GEN_43 = T_1525;
  assign GEN_413 = write ? GEN_43 : enables_0_6;
  assign T_1529 = masked_wdata[7];
  assign GEN_44 = T_1529;
  assign GEN_416 = write ? GEN_44 : enables_0_7;
  assign T_1533 = masked_wdata[8];
  assign GEN_45 = T_1533;
  assign GEN_419 = write ? GEN_45 : enables_0_8;
  assign T_1537 = masked_wdata[9];
  assign GEN_46 = T_1537;
  assign GEN_422 = write ? GEN_46 : enables_0_9;
  assign T_1541 = masked_wdata[10];
  assign GEN_47 = T_1541;
  assign GEN_425 = write ? GEN_47 : enables_0_10;
  assign T_1545 = masked_wdata[11];
  assign GEN_48 = T_1545;
  assign GEN_428 = write ? GEN_48 : enables_0_11;
  assign T_1549 = masked_wdata[12];
  assign GEN_49 = T_1549;
  assign GEN_431 = write ? GEN_49 : enables_0_12;
  assign T_1553 = masked_wdata[13];
  assign GEN_50 = T_1553;
  assign GEN_434 = write ? GEN_50 : enables_0_13;
  assign T_1557 = masked_wdata[14];
  assign GEN_51 = T_1557;
  assign GEN_437 = write ? GEN_51 : enables_0_14;
  assign T_1561 = masked_wdata[15];
  assign GEN_52 = T_1561;
  assign GEN_440 = write ? GEN_52 : enables_0_15;
  assign T_1565 = masked_wdata[16];
  assign GEN_53 = T_1565;
  assign GEN_443 = write ? GEN_53 : enables_0_16;
  assign T_1569 = masked_wdata[17];
  assign GEN_54 = T_1569;
  assign GEN_446 = write ? GEN_54 : enables_0_17;
  assign T_1573 = masked_wdata[18];
  assign GEN_55 = T_1573;
  assign GEN_449 = write ? GEN_55 : enables_0_18;
  assign T_1577 = masked_wdata[19];
  assign GEN_56 = T_1577;
  assign GEN_452 = write ? GEN_56 : enables_0_19;
  assign T_1581 = masked_wdata[20];
  assign GEN_57 = T_1581;
  assign GEN_455 = write ? GEN_57 : enables_0_20;
  assign T_1585 = masked_wdata[21];
  assign GEN_58 = T_1585;
  assign GEN_458 = write ? GEN_58 : enables_0_21;
  assign T_1589 = masked_wdata[22];
  assign GEN_59 = T_1589;
  assign GEN_461 = write ? GEN_59 : enables_0_22;
  assign T_1593 = masked_wdata[23];
  assign GEN_60 = T_1593;
  assign GEN_464 = write ? GEN_60 : enables_0_23;
  assign T_1597 = masked_wdata[24];
  assign GEN_61 = T_1597;
  assign GEN_467 = write ? GEN_61 : enables_0_24;
  assign T_1601 = masked_wdata[25];
  assign GEN_62 = T_1601;
  assign GEN_470 = write ? GEN_62 : enables_0_25;
  assign T_1605 = masked_wdata[26];
  assign GEN_63 = T_1605;
  assign GEN_473 = write ? GEN_63 : enables_0_26;
  assign T_1609 = masked_wdata[27];
  assign GEN_64 = T_1609;
  assign GEN_476 = write ? GEN_64 : enables_0_27;
  assign T_1613 = masked_wdata[28];
  assign GEN_65 = T_1613;
  assign GEN_479 = write ? GEN_65 : enables_0_28;
  assign T_1617 = masked_wdata[29];
  assign GEN_66 = T_1617;
  assign GEN_482 = write ? GEN_66 : enables_0_29;
  assign T_1621 = masked_wdata[30];
  assign GEN_67 = T_1621;
  assign GEN_485 = write ? GEN_67 : enables_0_30;
  assign T_1625 = masked_wdata[31];
  assign GEN_68 = T_1625;
  assign GEN_488 = write ? GEN_68 : enables_0_31;
  assign GEN_521 = {{32'd0}, T_1497};
  assign GEN_619 = T_1462 ? GEN_521 : GEN_326;
  assign GEN_623 = T_1462 ? GEN_398 : enables_0_1;
  assign GEN_625 = T_1462 ? GEN_401 : enables_0_2;
  assign GEN_627 = T_1462 ? GEN_404 : enables_0_3;
  assign GEN_629 = T_1462 ? GEN_407 : enables_0_4;
  assign GEN_631 = T_1462 ? GEN_410 : enables_0_5;
  assign GEN_633 = T_1462 ? GEN_413 : enables_0_6;
  assign GEN_635 = T_1462 ? GEN_416 : enables_0_7;
  assign GEN_637 = T_1462 ? GEN_419 : enables_0_8;
  assign GEN_639 = T_1462 ? GEN_422 : enables_0_9;
  assign GEN_641 = T_1462 ? GEN_425 : enables_0_10;
  assign GEN_643 = T_1462 ? GEN_428 : enables_0_11;
  assign GEN_645 = T_1462 ? GEN_431 : enables_0_12;
  assign GEN_647 = T_1462 ? GEN_434 : enables_0_13;
  assign GEN_649 = T_1462 ? GEN_437 : enables_0_14;
  assign GEN_651 = T_1462 ? GEN_440 : enables_0_15;
  assign GEN_653 = T_1462 ? GEN_443 : enables_0_16;
  assign GEN_655 = T_1462 ? GEN_446 : enables_0_17;
  assign GEN_657 = T_1462 ? GEN_449 : enables_0_18;
  assign GEN_659 = T_1462 ? GEN_452 : enables_0_19;
  assign GEN_661 = T_1462 ? GEN_455 : enables_0_20;
  assign GEN_663 = T_1462 ? GEN_458 : enables_0_21;
  assign GEN_665 = T_1462 ? GEN_461 : enables_0_22;
  assign GEN_667 = T_1462 ? GEN_464 : enables_0_23;
  assign GEN_669 = T_1462 ? GEN_467 : enables_0_24;
  assign GEN_671 = T_1462 ? GEN_470 : enables_0_25;
  assign GEN_673 = T_1462 ? GEN_473 : enables_0_26;
  assign GEN_675 = T_1462 ? GEN_476 : enables_0_27;
  assign GEN_677 = T_1462 ? GEN_479 : enables_0_28;
  assign GEN_679 = T_1462 ? GEN_482 : enables_0_29;
  assign GEN_681 = T_1462 ? GEN_485 : enables_0_30;
  assign GEN_683 = T_1462 ? GEN_488 : enables_0_31;
  assign T_1627 = addr >= 26'h1000;
  assign T_1631 = T_1459 == 1'h0;
  assign T_1632 = T_1461 & T_1631;
  assign T_1633 = T_1632 & T_1627;
  assign T_1634 = addr[4:3];
  assign T_1635 = {pending_1,pending_0};
  assign T_1636 = {pending_3,pending_2};
  assign T_1637 = {T_1636,T_1635};
  assign T_1638 = {pending_5,pending_4};
  assign T_1639 = {pending_7,pending_6};
  assign T_1640 = {T_1639,T_1638};
  assign T_1641 = {T_1640,T_1637};
  assign T_1642 = {pending_9,pending_8};
  assign T_1643 = {pending_11,pending_10};
  assign T_1644 = {T_1643,T_1642};
  assign T_1645 = {pending_13,pending_12};
  assign T_1646 = {pending_15,pending_14};
  assign T_1647 = {T_1646,T_1645};
  assign T_1648 = {T_1647,T_1644};
  assign T_1649 = {T_1648,T_1641};
  assign T_1650 = {pending_17,pending_16};
  assign T_1651 = {pending_19,pending_18};
  assign T_1652 = {T_1651,T_1650};
  assign T_1653 = {pending_21,pending_20};
  assign T_1654 = {pending_23,pending_22};
  assign T_1655 = {T_1654,T_1653};
  assign T_1656 = {T_1655,T_1652};
  assign T_1657 = {pending_25,pending_24};
  assign T_1658 = {pending_27,pending_26};
  assign T_1659 = {T_1658,T_1657};
  assign T_1660 = {pending_29,pending_28};
  assign T_1661 = {pending_31,pending_30};
  assign T_1662 = {T_1661,T_1660};
  assign T_1663 = {T_1662,T_1659};
  assign T_1664 = {T_1663,T_1656};
  assign T_1665 = {T_1664,T_1649};
  assign GEN_779 = {{5'd0}, T_1634};
  assign T_1667 = GEN_779 * 7'h40;
  assign T_1668 = T_1665 >> T_1667;
  assign GEN_684 = T_1633 ? {{32'd0}, T_1668} : GEN_619;
  assign T_1675 = T_1627 == 1'h0;
  assign T_1676 = T_1632 & T_1675;
  assign T_1677 = addr[6:3];
  assign T_1679 = T_1677 == 4'h0;
  assign T_1681 = {31'h0,priority_0};
  assign T_1683 = {31'h0,priority_1};
  assign T_1684 = {T_1683,T_1681};
  assign GEN_685 = T_1679 ? T_1684 : GEN_684;
  assign T_1686 = T_1677 == 4'h1;
  assign T_1688 = {31'h0,priority_2};
  assign T_1690 = {31'h0,priority_3};
  assign T_1691 = {T_1690,T_1688};
  assign GEN_686 = T_1686 ? T_1691 : GEN_685;
  assign T_1693 = T_1677 == 4'h2;
  assign T_1695 = {31'h0,priority_4};
  assign T_1697 = {31'h0,priority_5};
  assign T_1698 = {T_1697,T_1695};
  assign GEN_687 = T_1693 ? T_1698 : GEN_686;
  assign T_1700 = T_1677 == 4'h3;
  assign T_1702 = {31'h0,priority_6};
  assign T_1704 = {31'h0,priority_7};
  assign T_1705 = {T_1704,T_1702};
  assign GEN_688 = T_1700 ? T_1705 : GEN_687;
  assign T_1707 = T_1677 == 4'h4;
  assign T_1709 = {31'h0,priority_8};
  assign T_1711 = {31'h0,priority_9};
  assign T_1712 = {T_1711,T_1709};
  assign GEN_689 = T_1707 ? T_1712 : GEN_688;
  assign T_1714 = T_1677 == 4'h5;
  assign T_1716 = {31'h0,priority_10};
  assign T_1718 = {31'h0,priority_11};
  assign T_1719 = {T_1718,T_1716};
  assign GEN_690 = T_1714 ? T_1719 : GEN_689;
  assign T_1721 = T_1677 == 4'h6;
  assign T_1723 = {31'h0,priority_12};
  assign T_1725 = {31'h0,priority_13};
  assign T_1726 = {T_1725,T_1723};
  assign GEN_691 = T_1721 ? T_1726 : GEN_690;
  assign T_1728 = T_1677 == 4'h7;
  assign T_1730 = {31'h0,priority_14};
  assign T_1732 = {31'h0,priority_15};
  assign T_1733 = {T_1732,T_1730};
  assign GEN_692 = T_1728 ? T_1733 : GEN_691;
  assign T_1735 = T_1677 == 4'h8;
  assign T_1737 = {31'h0,priority_16};
  assign T_1739 = {31'h0,priority_17};
  assign T_1740 = {T_1739,T_1737};
  assign GEN_693 = T_1735 ? T_1740 : GEN_692;
  assign T_1742 = T_1677 == 4'h9;
  assign T_1744 = {31'h0,priority_18};
  assign T_1746 = {31'h0,priority_19};
  assign T_1747 = {T_1746,T_1744};
  assign GEN_694 = T_1742 ? T_1747 : GEN_693;
  assign T_1749 = T_1677 == 4'ha;
  assign T_1751 = {31'h0,priority_20};
  assign T_1753 = {31'h0,priority_21};
  assign T_1754 = {T_1753,T_1751};
  assign GEN_695 = T_1749 ? T_1754 : GEN_694;
  assign T_1756 = T_1677 == 4'hb;
  assign T_1758 = {31'h0,priority_22};
  assign T_1760 = {31'h0,priority_23};
  assign T_1761 = {T_1760,T_1758};
  assign GEN_696 = T_1756 ? T_1761 : GEN_695;
  assign T_1763 = T_1677 == 4'hc;
  assign T_1765 = {31'h0,priority_24};
  assign T_1767 = {31'h0,priority_25};
  assign T_1768 = {T_1767,T_1765};
  assign GEN_697 = T_1763 ? T_1768 : GEN_696;
  assign T_1770 = T_1677 == 4'hd;
  assign T_1772 = {31'h0,priority_26};
  assign T_1774 = {31'h0,priority_27};
  assign T_1775 = {T_1774,T_1772};
  assign GEN_698 = T_1770 ? T_1775 : GEN_697;
  assign T_1777 = T_1677 == 4'he;
  assign T_1779 = {31'h0,priority_28};
  assign T_1781 = {31'h0,priority_29};
  assign T_1782 = {T_1781,T_1779};
  assign GEN_699 = T_1777 ? T_1782 : GEN_698;
  assign T_1784 = T_1677 == 4'hf;
  assign T_1786 = {31'h0,priority_30};
  assign T_1788 = {31'h0,priority_31};
  assign T_1789 = {T_1788,T_1786};
  assign GEN_700 = T_1784 ? T_1789 : GEN_699;
  assign GEN_701 = T_1676 ? GEN_700 : GEN_684;
  assign T_1809 = 3'h6 == acq_io_deq_bits_a_type;
  assign T_1810 = T_1809 ? 3'h1 : 3'h3;
  assign T_1811 = 3'h5 == acq_io_deq_bits_a_type;
  assign T_1812 = T_1811 ? 3'h1 : T_1810;
  assign T_1813 = 3'h4 == acq_io_deq_bits_a_type;
  assign T_1814 = T_1813 ? 3'h4 : T_1812;
  assign T_1815 = 3'h3 == acq_io_deq_bits_a_type;
  assign T_1816 = T_1815 ? 3'h3 : T_1814;
  assign T_1817 = 3'h2 == acq_io_deq_bits_a_type;
  assign T_1818 = T_1817 ? 3'h3 : T_1816;
  assign T_1819 = 3'h1 == acq_io_deq_bits_a_type;
  assign T_1820 = T_1819 ? 3'h5 : T_1818;
  assign T_1821 = 3'h0 == acq_io_deq_bits_a_type;
  assign T_1822 = T_1821 ? 3'h4 : T_1820;
  assign T_1847_addr_beat = 3'h0;
  assign T_1847_client_xact_id = acq_io_deq_bits_client_xact_id;
  assign T_1847_manager_xact_id = 1'h0;
  assign T_1847_is_builtin_type = 1'h1;
  assign T_1847_g_type = {{1'd0}, T_1822};
  assign T_1847_data = rdata;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_100 = {1{$random}};
  pending_0 = GEN_100[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_132 = {1{$random}};
  pending_1 = GEN_132[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_133 = {1{$random}};
  pending_2 = GEN_133[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_227 = {1{$random}};
  pending_3 = GEN_227[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_259 = {1{$random}};
  pending_4 = GEN_259[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_260 = {1{$random}};
  pending_5 = GEN_260[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_292 = {1{$random}};
  pending_6 = GEN_292[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_293 = {1{$random}};
  pending_7 = GEN_293[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_325 = {1{$random}};
  pending_8 = GEN_325[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_327 = {1{$random}};
  pending_9 = GEN_327[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_328 = {1{$random}};
  pending_10 = GEN_328[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_360 = {1{$random}};
  pending_11 = GEN_360[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_361 = {1{$random}};
  pending_12 = GEN_361[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_393 = {1{$random}};
  pending_13 = GEN_393[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_394 = {1{$random}};
  pending_14 = GEN_394[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_395 = {1{$random}};
  pending_15 = GEN_395[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_396 = {1{$random}};
  pending_16 = GEN_396[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_397 = {1{$random}};
  pending_17 = GEN_397[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_399 = {1{$random}};
  pending_18 = GEN_399[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_400 = {1{$random}};
  pending_19 = GEN_400[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_402 = {1{$random}};
  pending_20 = GEN_402[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_403 = {1{$random}};
  pending_21 = GEN_403[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_405 = {1{$random}};
  pending_22 = GEN_405[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_406 = {1{$random}};
  pending_23 = GEN_406[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_408 = {1{$random}};
  pending_24 = GEN_408[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_409 = {1{$random}};
  pending_25 = GEN_409[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_411 = {1{$random}};
  pending_26 = GEN_411[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_412 = {1{$random}};
  pending_27 = GEN_412[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_414 = {1{$random}};
  pending_28 = GEN_414[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_415 = {1{$random}};
  pending_29 = GEN_415[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_417 = {1{$random}};
  pending_30 = GEN_417[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_418 = {1{$random}};
  pending_31 = GEN_418[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_420 = {1{$random}};
  enables_0_0 = GEN_420[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_421 = {1{$random}};
  enables_0_1 = GEN_421[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_423 = {1{$random}};
  enables_0_2 = GEN_423[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_424 = {1{$random}};
  enables_0_3 = GEN_424[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_426 = {1{$random}};
  enables_0_4 = GEN_426[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_427 = {1{$random}};
  enables_0_5 = GEN_427[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_429 = {1{$random}};
  enables_0_6 = GEN_429[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_430 = {1{$random}};
  enables_0_7 = GEN_430[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_432 = {1{$random}};
  enables_0_8 = GEN_432[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_433 = {1{$random}};
  enables_0_9 = GEN_433[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_435 = {1{$random}};
  enables_0_10 = GEN_435[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_436 = {1{$random}};
  enables_0_11 = GEN_436[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_438 = {1{$random}};
  enables_0_12 = GEN_438[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_439 = {1{$random}};
  enables_0_13 = GEN_439[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_441 = {1{$random}};
  enables_0_14 = GEN_441[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_442 = {1{$random}};
  enables_0_15 = GEN_442[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_444 = {1{$random}};
  enables_0_16 = GEN_444[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_445 = {1{$random}};
  enables_0_17 = GEN_445[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_447 = {1{$random}};
  enables_0_18 = GEN_447[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_448 = {1{$random}};
  enables_0_19 = GEN_448[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_450 = {1{$random}};
  enables_0_20 = GEN_450[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_451 = {1{$random}};
  enables_0_21 = GEN_451[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_453 = {1{$random}};
  enables_0_22 = GEN_453[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_454 = {1{$random}};
  enables_0_23 = GEN_454[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_456 = {1{$random}};
  enables_0_24 = GEN_456[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_457 = {1{$random}};
  enables_0_25 = GEN_457[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_459 = {1{$random}};
  enables_0_26 = GEN_459[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_460 = {1{$random}};
  enables_0_27 = GEN_460[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_462 = {1{$random}};
  enables_0_28 = GEN_462[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_463 = {1{$random}};
  enables_0_29 = GEN_463[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_465 = {1{$random}};
  enables_0_30 = GEN_465[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_466 = {1{$random}};
  enables_0_31 = GEN_466[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_468 = {1{$random}};
  T_1182 = GEN_468[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_469 = {1{$random}};
  T_1183 = GEN_469[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      pending_0 <= T_733_0;
    end else begin
      pending_0 <= 1'h0;
    end
    if(reset) begin
      pending_1 <= T_733_1;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h1 == myMaxDev) begin
            pending_1 <= GEN_2;
          end else begin
            if(io_devices_0_valid) begin
              pending_1 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_0_valid) begin
            pending_1 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_0_valid) begin
          pending_1 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_2 <= T_733_2;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h2 == myMaxDev) begin
            pending_2 <= GEN_2;
          end else begin
            if(io_devices_1_valid) begin
              pending_2 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_1_valid) begin
            pending_2 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_1_valid) begin
          pending_2 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_3 <= T_733_3;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h3 == myMaxDev) begin
            pending_3 <= GEN_2;
          end else begin
            if(io_devices_2_valid) begin
              pending_3 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_2_valid) begin
            pending_3 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_2_valid) begin
          pending_3 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_4 <= T_733_4;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h4 == myMaxDev) begin
            pending_4 <= GEN_2;
          end else begin
            if(io_devices_3_valid) begin
              pending_4 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_3_valid) begin
            pending_4 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_3_valid) begin
          pending_4 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_5 <= T_733_5;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h5 == myMaxDev) begin
            pending_5 <= GEN_2;
          end else begin
            if(io_devices_4_valid) begin
              pending_5 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_4_valid) begin
            pending_5 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_4_valid) begin
          pending_5 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_6 <= T_733_6;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h6 == myMaxDev) begin
            pending_6 <= GEN_2;
          end else begin
            if(io_devices_5_valid) begin
              pending_6 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_5_valid) begin
            pending_6 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_5_valid) begin
          pending_6 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_7 <= T_733_7;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h7 == myMaxDev) begin
            pending_7 <= GEN_2;
          end else begin
            if(io_devices_6_valid) begin
              pending_7 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_6_valid) begin
            pending_7 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_6_valid) begin
          pending_7 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_8 <= T_733_8;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h8 == myMaxDev) begin
            pending_8 <= GEN_2;
          end else begin
            if(io_devices_7_valid) begin
              pending_8 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_7_valid) begin
            pending_8 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_7_valid) begin
          pending_8 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_9 <= T_733_9;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h9 == myMaxDev) begin
            pending_9 <= GEN_2;
          end else begin
            if(io_devices_8_valid) begin
              pending_9 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_8_valid) begin
            pending_9 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_8_valid) begin
          pending_9 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_10 <= T_733_10;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'ha == myMaxDev) begin
            pending_10 <= GEN_2;
          end else begin
            if(io_devices_9_valid) begin
              pending_10 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_9_valid) begin
            pending_10 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_9_valid) begin
          pending_10 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_11 <= T_733_11;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'hb == myMaxDev) begin
            pending_11 <= GEN_2;
          end else begin
            if(io_devices_10_valid) begin
              pending_11 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_10_valid) begin
            pending_11 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_10_valid) begin
          pending_11 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_12 <= T_733_12;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'hc == myMaxDev) begin
            pending_12 <= GEN_2;
          end else begin
            if(io_devices_11_valid) begin
              pending_12 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_11_valid) begin
            pending_12 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_11_valid) begin
          pending_12 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_13 <= T_733_13;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'hd == myMaxDev) begin
            pending_13 <= GEN_2;
          end else begin
            if(io_devices_12_valid) begin
              pending_13 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_12_valid) begin
            pending_13 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_12_valid) begin
          pending_13 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_14 <= T_733_14;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'he == myMaxDev) begin
            pending_14 <= GEN_2;
          end else begin
            if(io_devices_13_valid) begin
              pending_14 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_13_valid) begin
            pending_14 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_13_valid) begin
          pending_14 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_15 <= T_733_15;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'hf == myMaxDev) begin
            pending_15 <= GEN_2;
          end else begin
            if(io_devices_14_valid) begin
              pending_15 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_14_valid) begin
            pending_15 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_14_valid) begin
          pending_15 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_16 <= T_733_16;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h10 == myMaxDev) begin
            pending_16 <= GEN_2;
          end else begin
            if(io_devices_15_valid) begin
              pending_16 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_15_valid) begin
            pending_16 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_15_valid) begin
          pending_16 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_17 <= T_733_17;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h11 == myMaxDev) begin
            pending_17 <= GEN_2;
          end else begin
            if(io_devices_16_valid) begin
              pending_17 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_16_valid) begin
            pending_17 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_16_valid) begin
          pending_17 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_18 <= T_733_18;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h12 == myMaxDev) begin
            pending_18 <= GEN_2;
          end else begin
            if(io_devices_17_valid) begin
              pending_18 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_17_valid) begin
            pending_18 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_17_valid) begin
          pending_18 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_19 <= T_733_19;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h13 == myMaxDev) begin
            pending_19 <= GEN_2;
          end else begin
            if(io_devices_18_valid) begin
              pending_19 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_18_valid) begin
            pending_19 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_18_valid) begin
          pending_19 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_20 <= T_733_20;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h14 == myMaxDev) begin
            pending_20 <= GEN_2;
          end else begin
            if(io_devices_19_valid) begin
              pending_20 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_19_valid) begin
            pending_20 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_19_valid) begin
          pending_20 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_21 <= T_733_21;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h15 == myMaxDev) begin
            pending_21 <= GEN_2;
          end else begin
            if(io_devices_20_valid) begin
              pending_21 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_20_valid) begin
            pending_21 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_20_valid) begin
          pending_21 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_22 <= T_733_22;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h16 == myMaxDev) begin
            pending_22 <= GEN_2;
          end else begin
            if(io_devices_21_valid) begin
              pending_22 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_21_valid) begin
            pending_22 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_21_valid) begin
          pending_22 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_23 <= T_733_23;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h17 == myMaxDev) begin
            pending_23 <= GEN_2;
          end else begin
            if(io_devices_22_valid) begin
              pending_23 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_22_valid) begin
            pending_23 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_22_valid) begin
          pending_23 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_24 <= T_733_24;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h18 == myMaxDev) begin
            pending_24 <= GEN_2;
          end else begin
            if(io_devices_23_valid) begin
              pending_24 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_23_valid) begin
            pending_24 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_23_valid) begin
          pending_24 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_25 <= T_733_25;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h19 == myMaxDev) begin
            pending_25 <= GEN_2;
          end else begin
            if(io_devices_24_valid) begin
              pending_25 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_24_valid) begin
            pending_25 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_24_valid) begin
          pending_25 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_26 <= T_733_26;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h1a == myMaxDev) begin
            pending_26 <= GEN_2;
          end else begin
            if(io_devices_25_valid) begin
              pending_26 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_25_valid) begin
            pending_26 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_25_valid) begin
          pending_26 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_27 <= T_733_27;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h1b == myMaxDev) begin
            pending_27 <= GEN_2;
          end else begin
            if(io_devices_26_valid) begin
              pending_27 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_26_valid) begin
            pending_27 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_26_valid) begin
          pending_27 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_28 <= T_733_28;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h1c == myMaxDev) begin
            pending_28 <= GEN_2;
          end else begin
            if(io_devices_27_valid) begin
              pending_28 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_27_valid) begin
            pending_28 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_27_valid) begin
          pending_28 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_29 <= T_733_29;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h1d == myMaxDev) begin
            pending_29 <= GEN_2;
          end else begin
            if(io_devices_28_valid) begin
              pending_29 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_28_valid) begin
            pending_29 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_28_valid) begin
          pending_29 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_30 <= T_733_30;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h1e == myMaxDev) begin
            pending_30 <= GEN_2;
          end else begin
            if(io_devices_29_valid) begin
              pending_30 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_29_valid) begin
            pending_30 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_29_valid) begin
          pending_30 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_31 <= T_733_31;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h1f == myMaxDev) begin
            pending_31 <= GEN_2;
          end else begin
            if(io_devices_30_valid) begin
              pending_31 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_30_valid) begin
            pending_31 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_30_valid) begin
          pending_31 <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      enables_0_0 <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_1 <= GEN_38;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_2 <= GEN_39;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_3 <= GEN_40;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_4 <= GEN_41;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_5 <= GEN_42;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_6 <= GEN_43;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_7 <= GEN_44;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_8 <= GEN_45;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_9 <= GEN_46;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_10 <= GEN_47;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_11 <= GEN_48;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_12 <= GEN_49;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_13 <= GEN_50;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_14 <= GEN_51;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_15 <= GEN_52;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_16 <= GEN_53;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_17 <= GEN_54;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_18 <= GEN_55;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_19 <= GEN_56;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_20 <= GEN_57;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_21 <= GEN_58;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_22 <= GEN_59;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_23 <= GEN_60;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_24 <= GEN_61;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_25 <= GEN_62;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_26 <= GEN_63;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_27 <= GEN_64;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_28 <= GEN_65;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_29 <= GEN_66;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_30 <= GEN_67;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_31 <= GEN_68;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1176) begin
        T_1182 <= {{1'd0}, T_1069};
      end else begin
        T_1182 <= T_1180;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1176) begin
        if(T_1064) begin
          if(T_1008) begin
            if(T_980) begin
              if(T_966) begin
                T_1183 <= 2'h2;
              end else begin
                T_1183 <= T_901;
              end
            end else begin
              if(T_974) begin
                T_1183 <= T_903;
              end else begin
                T_1183 <= T_905;
              end
            end
          end else begin
            if(T_1002) begin
              if(T_988) begin
                T_1183 <= T_907;
              end else begin
                T_1183 <= T_909;
              end
            end else begin
              if(T_996) begin
                T_1183 <= T_911;
              end else begin
                T_1183 <= T_913;
              end
            end
          end
        end else begin
          if(T_1058) begin
            if(T_1030) begin
              if(T_1016) begin
                T_1183 <= T_915;
              end else begin
                T_1183 <= T_917;
              end
            end else begin
              if(T_1024) begin
                T_1183 <= T_919;
              end else begin
                T_1183 <= T_921;
              end
            end
          end else begin
            if(T_1052) begin
              if(T_1038) begin
                T_1183 <= T_923;
              end else begin
                T_1183 <= T_925;
              end
            end else begin
              if(T_1046) begin
                T_1183 <= T_927;
              end else begin
                T_1183 <= T_929;
              end
            end
          end
        end
      end else begin
        if(T_1170) begin
          if(T_1114) begin
            if(T_1086) begin
              if(T_1072) begin
                T_1183 <= T_931;
              end else begin
                T_1183 <= T_933;
              end
            end else begin
              if(T_1080) begin
                T_1183 <= T_935;
              end else begin
                T_1183 <= T_937;
              end
            end
          end else begin
            if(T_1108) begin
              if(T_1094) begin
                T_1183 <= T_939;
              end else begin
                T_1183 <= T_941;
              end
            end else begin
              if(T_1102) begin
                T_1183 <= T_943;
              end else begin
                T_1183 <= T_945;
              end
            end
          end
        end else begin
          if(T_1164) begin
            if(T_1136) begin
              if(T_1122) begin
                T_1183 <= T_947;
              end else begin
                T_1183 <= T_949;
              end
            end else begin
              if(T_1130) begin
                T_1183 <= T_951;
              end else begin
                T_1183 <= T_953;
              end
            end
          end else begin
            if(T_1158) begin
              if(T_1144) begin
                T_1183 <= T_955;
              end else begin
                T_1183 <= T_957;
              end
            end else begin
              if(T_1152) begin
                T_1183 <= T_959;
              end else begin
                T_1183 <= T_961;
              end
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1225) begin
          $fwrite(32'h80000002,"Assertion failed: unsupported PLIC operation\n    at Plic.scala:108 assert(!acq.fire() || read || write, ---unsupported PLIC operation---)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module LevelGateway(
  input   clk,
  input   reset,
  input   io_interrupt,
  output  io_plic_valid,
  input   io_plic_ready,
  input   io_plic_complete
);
  reg  inFlight;
  reg [31:0] GEN_2;
  wire  T_6;
  wire  GEN_0;
  wire  GEN_1;
  wire  T_10;
  wire  T_11;
  assign io_plic_valid = T_11;
  assign T_6 = io_interrupt & io_plic_ready;
  assign GEN_0 = T_6 ? 1'h1 : inFlight;
  assign GEN_1 = io_plic_complete ? 1'h0 : GEN_0;
  assign T_10 = inFlight == 1'h0;
  assign T_11 = io_interrupt & T_10;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_2 = {1{$random}};
  inFlight = GEN_2[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      inFlight <= 1'h0;
    end else begin
      if(io_plic_complete) begin
        inFlight <= 1'h0;
      end else begin
        if(T_6) begin
          inFlight <= 1'h1;
        end
      end
    end
  end
endmodule
module DebugModule(
  input   clk,
  input   reset,
  output  io_db_req_ready,
  input   io_db_req_valid,
  input  [4:0] io_db_req_bits_addr,
  input  [1:0] io_db_req_bits_op,
  input  [33:0] io_db_req_bits_data,
  input   io_db_resp_ready,
  output  io_db_resp_valid,
  output [1:0] io_db_resp_bits_resp,
  output [33:0] io_db_resp_bits_data,
  output  io_debugInterrupts_0,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [11:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data,
  output  io_ndreset,
  output  io_fullreset
);
  wire  CONTROLReset_interrupt;
  wire  CONTROLReset_haltnot;
  wire [9:0] CONTROLReset_reserved0;
  wire [2:0] CONTROLReset_buserror;
  wire [2:0] CONTROLReset_serial;
  wire  CONTROLReset_autoincrement;
  wire [2:0] CONTROLReset_access;
  wire [9:0] CONTROLReset_hartid;
  wire  CONTROLReset_ndreset;
  wire  CONTROLReset_fullreset;
  wire  CONTROLWrEn;
  reg  CONTROLReg_interrupt;
  reg [31:0] GEN_26;
  reg  CONTROLReg_haltnot;
  reg [31:0] GEN_27;
  reg [9:0] CONTROLReg_reserved0;
  reg [31:0] GEN_28;
  reg [2:0] CONTROLReg_buserror;
  reg [31:0] GEN_29;
  reg [2:0] CONTROLReg_serial;
  reg [31:0] GEN_30;
  reg  CONTROLReg_autoincrement;
  reg [31:0] GEN_52;
  reg [2:0] CONTROLReg_access;
  reg [31:0] GEN_85;
  reg [9:0] CONTROLReg_hartid;
  reg [31:0] GEN_86;
  reg  CONTROLReg_ndreset;
  reg [31:0] GEN_88;
  reg  CONTROLReg_fullreset;
  reg [31:0] GEN_89;
  wire  CONTROLWrData_interrupt;
  wire  CONTROLWrData_haltnot;
  wire [9:0] CONTROLWrData_reserved0;
  wire [2:0] CONTROLWrData_buserror;
  wire [2:0] CONTROLWrData_serial;
  wire  CONTROLWrData_autoincrement;
  wire [2:0] CONTROLWrData_access;
  wire [9:0] CONTROLWrData_hartid;
  wire  CONTROLWrData_ndreset;
  wire  CONTROLWrData_fullreset;
  wire  CONTROLRdData_interrupt;
  wire  CONTROLRdData_haltnot;
  wire [9:0] CONTROLRdData_reserved0;
  wire [2:0] CONTROLRdData_buserror;
  wire [2:0] CONTROLRdData_serial;
  wire  CONTROLRdData_autoincrement;
  wire [2:0] CONTROLRdData_access;
  wire [9:0] CONTROLRdData_hartid;
  wire  CONTROLRdData_ndreset;
  wire  CONTROLRdData_fullreset;
  reg  ndresetCtrReg;
  reg [31:0] GEN_90;
  wire [1:0] DMINFORdData_reserved0;
  wire [6:0] DMINFORdData_abussize;
  wire [3:0] DMINFORdData_serialcount;
  wire  DMINFORdData_access128;
  wire  DMINFORdData_access64;
  wire  DMINFORdData_access32;
  wire  DMINFORdData_access16;
  wire  DMINFORdData_accesss8;
  wire [5:0] DMINFORdData_dramsize;
  wire  DMINFORdData_haltsum;
  wire [2:0] DMINFORdData_reserved1;
  wire  DMINFORdData_authenticated;
  wire  DMINFORdData_authbusy;
  wire [1:0] DMINFORdData_authtype;
  wire [1:0] DMINFORdData_version;
  wire  HALTSUMRdData_serialfull;
  wire  HALTSUMRdData_serialvalid;
  wire [31:0] HALTSUMRdData_acks;
  wire  RAMWrData_interrupt;
  wire  RAMWrData_haltnot;
  wire [31:0] RAMWrData_data;
  wire  RAMRdData_interrupt;
  wire  RAMRdData_haltnot;
  wire [31:0] RAMRdData_data;
  wire  SETHALTNOTWrEn;
  wire [9:0] SETHALTNOTWrData;
  wire  CLEARDEBINTWrEn;
  wire [9:0] CLEARDEBINTWrData;
  wire  T_655_0;
  reg  interruptRegs_0;
  reg [31:0] GEN_109;
  wire  T_666_0;
  reg  haltnotRegs_0;
  reg [31:0] GEN_110;
  wire [31:0] haltnotStatus_0;
  wire [31:0] rdHaltnotStatus;
  wire  haltnotSummary;
  reg [63:0] ramMem [0:3];
  reg [63:0] GEN_111;
  wire [63:0] ramMem_T_850_data;
  wire [1:0] ramMem_T_850_addr;
  wire  ramMem_T_850_en;
  wire [63:0] ramMem_T_851_data;
  wire [1:0] ramMem_T_851_addr;
  wire  ramMem_T_851_mask;
  wire  ramMem_T_851_en;
  wire [1:0] ramAddr;
  wire [63:0] ramRdData;
  wire [63:0] ramWrData;
  wire [63:0] ramWrMask;
  wire  ramWrEn;
  wire [2:0] dbRamAddr;
  wire [31:0] dbRamRdData;
  wire [31:0] dbRamWrData;
  wire  dbRamWrEn;
  wire  dbRamRdEn;
  wire [1:0] sbRamAddr;
  wire [63:0] sbRamRdData;
  wire [63:0] sbRamWrData;
  wire  sbRamWrEn;
  wire  sbRamRdEn;
  wire [63:0] sbRomRdData;
  wire  dbRdEn;
  wire  dbWrEn;
  wire [33:0] dbRdData;
  reg  dbStateReg;
  reg [31:0] GEN_112;
  wire [1:0] dbResult_resp;
  wire [33:0] dbResult_data;
  wire [4:0] dbReq_addr;
  wire [1:0] dbReq_op;
  wire [33:0] dbReq_data;
  reg [1:0] dbRespReg_resp;
  reg [31:0] GEN_113;
  reg [33:0] dbRespReg_data;
  reg [63:0] GEN_114;
  wire  rdCondWrFailure;
  wire  dbWrNeeded;
  wire [11:0] sbAddr;
  wire [63:0] sbRdData;
  wire [63:0] sbWrData;
  wire [63:0] sbWrMask;
  wire  sbWrEn;
  wire  sbRdEn;
  wire  stallFromDb;
  wire  stallFromSb;
  wire  T_720;
  wire  T_721;
  wire  GEN_11;
  wire  GEN_12;
  wire  T_723;
  wire  T_724;
  wire  T_726;
  wire  T_727;
  wire  GEN_13;
  wire  GEN_14;
  wire  T_731;
  wire  T_732;
  wire  T_733;
  wire  T_735;
  wire  GEN_15;
  wire  GEN_16;
  wire  T_738;
  wire  GEN_17;
  wire  GEN_18;
  wire  T_741;
  wire  T_742;
  wire  T_745;
  wire  GEN_19;
  wire  GEN_20;
  wire  T_750;
  wire  T_751;
  wire  T_754;
  wire  GEN_21;
  wire  GEN_22;
  wire [2:0] T_782;
  wire [1:0] T_783;
  wire [31:0] T_799_0;
  wire [31:0] T_799_1;
  wire [31:0] dbRamWrMask_0;
  wire [31:0] dbRamWrMask_1;
  wire  T_804;
  wire [31:0] T_805;
  wire [31:0] T_806;
  wire [31:0] T_812_0;
  wire [31:0] T_812_1;
  wire [31:0] T_821_0;
  wire [31:0] T_821_1;
  wire [31:0] GEN_0;
  wire [31:0] GEN_23;
  wire [31:0] GEN_24;
  wire [31:0] GEN_1;
  wire [31:0] GEN_25;
  wire [63:0] T_828;
  wire [63:0] T_829;
  wire  T_830;
  wire  T_831;
  wire  T_832;
  wire  T_834;
  wire  T_835;
  wire  T_837;
  wire [63:0] dbRamWrDataVec;
  wire [63:0] T_838;
  wire [63:0] T_839;
  wire [63:0] T_840;
  wire [63:0] T_841;
  wire [63:0] T_842;
  wire [63:0] T_845;
  wire [63:0] T_846;
  wire  T_847;
  wire [1:0] T_848;
  wire [1:0] T_849;
  wire  T_852;
  wire  T_875_interrupt;
  wire  T_875_haltnot;
  wire [9:0] T_875_reserved0;
  wire [2:0] T_875_buserror;
  wire [2:0] T_875_serial;
  wire  T_875_autoincrement;
  wire [2:0] T_875_access;
  wire [9:0] T_875_hartid;
  wire  T_875_ndreset;
  wire  T_875_fullreset;
  wire  T_886;
  wire  T_887;
  wire [9:0] T_888;
  wire [2:0] T_889;
  wire  T_890;
  wire [2:0] T_891;
  wire [2:0] T_892;
  wire [9:0] T_893;
  wire  T_894;
  wire  T_895;
  wire  T_904_interrupt;
  wire  T_904_haltnot;
  wire [31:0] T_904_data;
  wire [31:0] T_908;
  wire  T_913;
  wire  T_915;
  wire  GEN_31;
  wire  T_917;
  wire  T_919;
  wire  T_920;
  wire  GEN_32;
  wire  T_924;
  wire  T_925;
  wire  GEN_33;
  wire  GEN_34;
  wire [9:0] GEN_35;
  wire [2:0] GEN_36;
  wire [2:0] GEN_37;
  wire  GEN_38;
  wire [2:0] GEN_39;
  wire [9:0] GEN_40;
  wire  GEN_41;
  wire  GEN_42;
  wire  GEN_43;
  wire  T_928;
  wire  T_929;
  wire  T_930;
  wire  GEN_44;
  wire  T_933;
  wire  T_935;
  wire [1:0] T_938;
  wire  T_939;
  wire  T_940;
  wire  GEN_45;
  wire [9:0] GEN_46;
  wire  GEN_47;
  wire  GEN_48;
  wire  T_945;
  wire  GEN_49;
  wire  GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire  T_958;
  wire [31:0] GEN_50;
  wire [1:0] T_963;
  wire [33:0] T_964;
  wire [33:0] GEN_51;
  wire [1:0] T_970;
  wire [3:0] T_971;
  wire [13:0] T_972;
  wire [15:0] T_973;
  wire [5:0] T_974;
  wire [1:0] T_975;
  wire [11:0] T_976;
  wire [17:0] T_977;
  wire [33:0] T_978;
  wire [33:0] GEN_53;
  wire  T_980;
  wire  T_986;
  wire [2:0] T_987;
  wire [4:0] T_988;
  wire [3:0] T_989;
  wire [6:0] T_990;
  wire [10:0] T_991;
  wire [15:0] T_992;
  wire [1:0] T_993;
  wire [1:0] T_994;
  wire [3:0] T_995;
  wire [4:0] T_996;
  wire [8:0] T_997;
  wire [13:0] T_998;
  wire [17:0] T_999;
  wire [33:0] T_1000;
  wire [33:0] GEN_54;
  wire  T_1002;
  wire  T_1009;
  wire  T_1010;
  wire  T_1011;
  wire [33:0] GEN_55;
  wire [2:0] T_1013;
  wire  T_1015;
  wire  T_1025;
  wire  T_1026;
  wire  T_1027;
  wire [33:0] GEN_56;
  wire  T_1040;
  wire  T_1041;
  wire [33:0] GEN_57;
  wire  T_1043;
  wire  T_1045;
  wire  T_1046;
  wire  T_1048;
  wire  T_1051;
  wire  T_1052;
  wire  T_1053;
  wire [1:0] T_1056;
  wire  T_1058;
  wire  T_1059;
  wire  T_1061;
  wire  T_1062;
  wire  T_1063;
  wire  T_1064;
  wire  T_1066;
  wire  T_1068;
  wire  GEN_58;
  wire [1:0] GEN_59;
  wire [33:0] GEN_60;
  wire  GEN_61;
  wire [1:0] GEN_62;
  wire [33:0] GEN_63;
  wire  T_1073;
  wire  T_1074;
  wire  GEN_64;
  wire [1:0] GEN_65;
  wire [33:0] GEN_66;
  wire  T_1078;
  wire  T_1079;
  wire  GEN_67;
  wire  GEN_68;
  wire [1:0] GEN_69;
  wire [33:0] GEN_70;
  wire [63:0] T_1101_0;
  wire [63:0] T_1101_1;
  wire [63:0] T_1101_2;
  wire [63:0] T_1101_3;
  wire [63:0] T_1101_4;
  wire [63:0] T_1101_5;
  wire [63:0] T_1101_6;
  wire [63:0] T_1101_7;
  wire [63:0] T_1101_8;
  wire [63:0] T_1101_9;
  wire [63:0] T_1101_10;
  wire [63:0] T_1101_11;
  wire [63:0] T_1101_12;
  wire [63:0] T_1101_13;
  wire [63:0] T_1101_14;
  wire [3:0] T_1104;
  wire [3:0] T_1105;
  wire [63:0] GEN_6;
  wire [63:0] GEN_71;
  wire [63:0] GEN_72;
  wire [63:0] GEN_73;
  wire [63:0] GEN_74;
  wire [63:0] GEN_75;
  wire [63:0] GEN_76;
  wire [63:0] GEN_77;
  wire [63:0] GEN_78;
  wire [63:0] GEN_79;
  wire [63:0] GEN_80;
  wire [63:0] GEN_81;
  wire [63:0] GEN_82;
  wire [63:0] GEN_83;
  wire [63:0] GEN_84;
  wire [31:0] T_1109;
  wire [31:0] T_1110;
  wire [31:0] T_1116_0;
  wire [31:0] T_1116_1;
  wire [31:0] T_1118;
  wire [31:0] T_1119;
  wire [31:0] T_1125_0;
  wire [31:0] T_1125_1;
  wire [31:0] GEN_7;
  wire [31:0] GEN_8;
  wire [3:0] T_1131;
  wire  T_1133;
  wire  GEN_87;
  wire [8:0] T_1134;
  wire  T_1137;
  wire [31:0] GEN_9;
  wire  T_1141;
  wire  T_1142;
  wire  T_1143;
  wire  T_1147;
  wire [31:0] GEN_10;
  wire  T_1151;
  wire  T_1152;
  wire  T_1153;
  wire [63:0] GEN_91;
  wire  GEN_92;
  wire  T_1162;
  wire  T_1165;
  wire  T_1166;
  wire  T_1168;
  wire  T_1169;
  wire [63:0] GEN_93;
  wire  T_1173;
  wire  T_1174;
  wire [63:0] GEN_94;
  reg [25:0] sbAcqReg_addr_block;
  reg [31:0] GEN_115;
  reg [1:0] sbAcqReg_client_xact_id;
  reg [31:0] GEN_116;
  reg [2:0] sbAcqReg_addr_beat;
  reg [31:0] GEN_117;
  reg  sbAcqReg_is_builtin_type;
  reg [31:0] GEN_118;
  reg [2:0] sbAcqReg_a_type;
  reg [31:0] GEN_119;
  reg [11:0] sbAcqReg_union;
  reg [31:0] GEN_120;
  reg [63:0] sbAcqReg_data;
  reg [63:0] GEN_121;
  reg  sbAcqValidReg;
  reg [31:0] GEN_122;
  wire  T_1203;
  wire  sbReg_get;
  wire  T_1204;
  wire  sbReg_getblk;
  wire  T_1205;
  wire  sbReg_put;
  wire  T_1206;
  wire  sbReg_putblk;
  wire  sbMultibeat;
  wire [3:0] T_1208;
  wire [2:0] sbBeatInc1;
  wire  sbLast;
  wire [2:0] T_1217_0;
  wire [2:0] T_1217_1;
  wire  T_1219;
  wire  T_1220;
  wire  T_1221;
  wire  T_1222;
  wire [2:0] T_1223;
  wire [2:0] T_1225;
  wire [28:0] T_1226;
  wire [31:0] T_1227;
  wire  T_1228;
  wire  T_1229;
  wire  T_1230;
  wire  T_1231;
  wire  T_1233;
  wire  T_1234;
  wire  T_1236;
  wire [1:0] T_1238;
  wire  T_1239;
  wire  T_1240;
  wire [3:0] T_1244;
  wire [3:0] T_1248;
  wire [7:0] T_1249;
  wire  T_1256;
  wire [7:0] T_1257;
  wire [7:0] T_1259;
  wire [7:0] T_1260;
  wire  T_1261;
  wire  T_1262;
  wire  T_1263;
  wire  T_1264;
  wire  T_1265;
  wire  T_1266;
  wire  T_1267;
  wire  T_1268;
  wire [7:0] T_1272;
  wire [7:0] T_1276;
  wire [7:0] T_1280;
  wire [7:0] T_1284;
  wire [7:0] T_1288;
  wire [7:0] T_1292;
  wire [7:0] T_1296;
  wire [7:0] T_1300;
  wire [15:0] T_1301;
  wire [15:0] T_1302;
  wire [31:0] T_1303;
  wire [15:0] T_1304;
  wire [15:0] T_1305;
  wire [31:0] T_1306;
  wire [63:0] T_1307;
  wire  T_1308;
  wire [25:0] GEN_95;
  wire [1:0] GEN_96;
  wire [2:0] GEN_97;
  wire  GEN_98;
  wire [2:0] GEN_99;
  wire [11:0] GEN_100;
  wire [63:0] GEN_101;
  wire  GEN_102;
  wire  T_1310;
  wire  T_1312;
  wire  T_1313;
  wire  GEN_103;
  wire [2:0] GEN_104;
  wire  GEN_105;
  wire  T_1316;
  wire  GEN_106;
  wire [2:0] GEN_107;
  wire  GEN_108;
  wire  T_1334;
  wire [2:0] T_1335;
  wire  T_1336;
  wire [2:0] T_1337;
  wire  T_1338;
  wire [2:0] T_1339;
  wire  T_1340;
  wire [2:0] T_1341;
  wire  T_1342;
  wire [2:0] T_1343;
  wire  T_1344;
  wire [2:0] T_1345;
  wire  T_1346;
  wire [2:0] T_1347;
  wire [2:0] T_1371_addr_beat;
  wire [1:0] T_1371_client_xact_id;
  wire  T_1371_manager_xact_id;
  wire  T_1371_is_builtin_type;
  wire [3:0] T_1371_g_type;
  wire [63:0] T_1371_data;
  wire  T_1396;
  wire  T_1397;
  wire  T_1399;
  wire  T_1400;
  wire  T_1401;
  wire  sbStall;
  wire  T_1403;
  assign io_db_req_ready = T_1064;
  assign io_db_resp_valid = dbStateReg;
  assign io_db_resp_bits_resp = dbRespReg_resp;
  assign io_db_resp_bits_data = dbRespReg_data;
  assign io_debugInterrupts_0 = interruptRegs_0;
  assign io_tl_acquire_ready = T_1403;
  assign io_tl_grant_valid = sbAcqValidReg;
  assign io_tl_grant_bits_addr_beat = T_1371_addr_beat;
  assign io_tl_grant_bits_client_xact_id = T_1371_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = T_1371_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = T_1371_is_builtin_type;
  assign io_tl_grant_bits_g_type = T_1371_g_type;
  assign io_tl_grant_bits_data = T_1371_data;
  assign io_ndreset = ndresetCtrReg;
  assign io_fullreset = CONTROLReg_fullreset;
  assign CONTROLReset_interrupt = 1'h0;
  assign CONTROLReset_haltnot = 1'h0;
  assign CONTROLReset_reserved0 = 10'h0;
  assign CONTROLReset_buserror = 3'h0;
  assign CONTROLReset_serial = 3'h0;
  assign CONTROLReset_autoincrement = 1'h0;
  assign CONTROLReset_access = 3'h2;
  assign CONTROLReset_hartid = 10'h0;
  assign CONTROLReset_ndreset = 1'h0;
  assign CONTROLReset_fullreset = 1'h0;
  assign CONTROLWrEn = GEN_32;
  assign CONTROLWrData_interrupt = T_875_interrupt;
  assign CONTROLWrData_haltnot = T_875_haltnot;
  assign CONTROLWrData_reserved0 = T_875_reserved0;
  assign CONTROLWrData_buserror = T_875_buserror;
  assign CONTROLWrData_serial = T_875_serial;
  assign CONTROLWrData_autoincrement = T_875_autoincrement;
  assign CONTROLWrData_access = T_875_access;
  assign CONTROLWrData_hartid = T_875_hartid;
  assign CONTROLWrData_ndreset = T_875_ndreset;
  assign CONTROLWrData_fullreset = T_875_fullreset;
  assign CONTROLRdData_interrupt = GEN_2;
  assign CONTROLRdData_haltnot = GEN_3;
  assign CONTROLRdData_reserved0 = CONTROLReg_reserved0;
  assign CONTROLRdData_buserror = CONTROLReg_buserror;
  assign CONTROLRdData_serial = CONTROLReg_serial;
  assign CONTROLRdData_autoincrement = CONTROLReg_autoincrement;
  assign CONTROLRdData_access = CONTROLReg_access;
  assign CONTROLRdData_hartid = CONTROLReg_hartid;
  assign CONTROLRdData_ndreset = ndresetCtrReg;
  assign CONTROLRdData_fullreset = CONTROLReg_fullreset;
  assign DMINFORdData_reserved0 = 2'h0;
  assign DMINFORdData_abussize = 7'h0;
  assign DMINFORdData_serialcount = 4'h0;
  assign DMINFORdData_access128 = 1'h0;
  assign DMINFORdData_access64 = 1'h0;
  assign DMINFORdData_access32 = 1'h0;
  assign DMINFORdData_access16 = 1'h0;
  assign DMINFORdData_accesss8 = 1'h0;
  assign DMINFORdData_dramsize = 6'h6;
  assign DMINFORdData_haltsum = 1'h0;
  assign DMINFORdData_reserved1 = 3'h0;
  assign DMINFORdData_authenticated = 1'h1;
  assign DMINFORdData_authbusy = 1'h0;
  assign DMINFORdData_authtype = 2'h0;
  assign DMINFORdData_version = 2'h1;
  assign HALTSUMRdData_serialfull = 1'h0;
  assign HALTSUMRdData_serialvalid = 1'h0;
  assign HALTSUMRdData_acks = {{31'd0}, haltnotSummary};
  assign RAMWrData_interrupt = T_904_interrupt;
  assign RAMWrData_haltnot = T_904_haltnot;
  assign RAMWrData_data = T_904_data;
  assign RAMRdData_interrupt = GEN_4;
  assign RAMRdData_haltnot = GEN_5;
  assign RAMRdData_data = dbRamRdData;
  assign SETHALTNOTWrEn = T_1143;
  assign SETHALTNOTWrData = GEN_7[9:0];
  assign CLEARDEBINTWrEn = T_1153;
  assign CLEARDEBINTWrData = GEN_8[9:0];
  assign T_655_0 = 1'h0;
  assign T_666_0 = 1'h0;
  assign haltnotStatus_0 = {{31'd0}, haltnotRegs_0};
  assign rdHaltnotStatus = GEN_50;
  assign haltnotSummary = haltnotStatus_0 != 32'h0;
  assign ramMem_T_850_addr = ramAddr;
  assign ramMem_T_850_en = 1'h1;
  assign ramMem_T_850_data = ramMem[ramMem_T_850_addr];
  assign ramMem_T_851_data = ramWrData;
  assign ramMem_T_851_addr = ramAddr;
  assign ramMem_T_851_mask = ramWrEn;
  assign ramMem_T_851_en = ramWrEn;
  assign ramAddr = T_849;
  assign ramRdData = ramMem_T_850_data;
  assign ramWrData = T_846;
  assign ramWrMask = T_829;
  assign ramWrEn = T_852;
  assign dbRamAddr = T_782;
  assign dbRamRdData = GEN_1;
  assign dbRamWrData = dbReq_data[31:0];
  assign dbRamWrEn = GEN_31;
  assign dbRamRdEn = 1'h0;
  assign sbRamAddr = T_783;
  assign sbRamRdData = ramRdData;
  assign sbRamWrData = sbWrData;
  assign sbRamWrEn = GEN_87;
  assign sbRamRdEn = GEN_92;
  assign sbRomRdData = GEN_6;
  assign dbRdEn = T_1066;
  assign dbWrEn = T_1068;
  assign dbRdData = GEN_57;
  assign dbResult_resp = T_1056;
  assign dbResult_data = dbRdData;
  assign dbReq_addr = io_db_req_bits_addr;
  assign dbReq_op = io_db_req_bits_op;
  assign dbReq_data = io_db_req_bits_data;
  assign rdCondWrFailure = T_1046;
  assign dbWrNeeded = T_1053;
  assign sbAddr = T_1227[11:0];
  assign sbRdData = GEN_94;
  assign sbWrData = sbAcqReg_data;
  assign sbWrMask = T_1307;
  assign sbWrEn = T_1231;
  assign sbRdEn = T_1229;
  assign stallFromDb = 1'h0;
  assign stallFromSb = T_831;
  assign T_720 = CONTROLWrData_hartid == 10'h0;
  assign T_721 = interruptRegs_0 | CONTROLWrData_interrupt;
  assign GEN_11 = T_720 ? T_721 : interruptRegs_0;
  assign GEN_12 = CONTROLWrEn ? GEN_11 : interruptRegs_0;
  assign T_723 = CONTROLWrEn == 1'h0;
  assign T_724 = T_723 & dbRamWrEn;
  assign T_726 = CONTROLReg_hartid == 10'h0;
  assign T_727 = interruptRegs_0 | RAMWrData_interrupt;
  assign GEN_13 = T_726 ? T_727 : GEN_12;
  assign GEN_14 = T_724 ? GEN_13 : GEN_12;
  assign T_731 = dbRamWrEn == 1'h0;
  assign T_732 = T_723 & T_731;
  assign T_733 = T_732 & CLEARDEBINTWrEn;
  assign T_735 = CLEARDEBINTWrData == 10'h0;
  assign GEN_15 = T_735 ? 1'h0 : GEN_14;
  assign GEN_16 = T_733 ? GEN_15 : GEN_14;
  assign T_738 = SETHALTNOTWrData == 10'h0;
  assign GEN_17 = T_738 ? 1'h1 : haltnotRegs_0;
  assign GEN_18 = SETHALTNOTWrEn ? GEN_17 : haltnotRegs_0;
  assign T_741 = SETHALTNOTWrEn == 1'h0;
  assign T_742 = T_741 & CONTROLWrEn;
  assign T_745 = haltnotRegs_0 & CONTROLWrData_haltnot;
  assign GEN_19 = T_720 ? T_745 : GEN_18;
  assign GEN_20 = T_742 ? GEN_19 : GEN_18;
  assign T_750 = T_741 & T_723;
  assign T_751 = T_750 & dbRamWrEn;
  assign T_754 = haltnotRegs_0 & RAMWrData_haltnot;
  assign GEN_21 = T_726 ? T_754 : GEN_20;
  assign GEN_22 = T_751 ? GEN_21 : GEN_20;
  assign T_782 = dbReq_addr[2:0];
  assign T_783 = sbAddr[4:3];
  assign T_799_0 = 32'hffffffff;
  assign T_799_1 = 32'hffffffff;
  assign dbRamWrMask_0 = GEN_23;
  assign dbRamWrMask_1 = GEN_24;
  assign T_804 = dbRamAddr[0];
  assign T_805 = ramRdData[31:0];
  assign T_806 = ramRdData[63:32];
  assign T_812_0 = T_805;
  assign T_812_1 = T_806;
  assign T_821_0 = 32'h0;
  assign T_821_1 = 32'h0;
  assign GEN_0 = 32'hffffffff;
  assign GEN_23 = 1'h0 == T_804 ? GEN_0 : T_821_0;
  assign GEN_24 = T_804 ? GEN_0 : T_821_1;
  assign GEN_1 = GEN_25;
  assign GEN_25 = T_804 ? T_812_1 : T_812_0;
  assign T_828 = {dbRamWrMask_1,dbRamWrMask_0};
  assign T_829 = sbRamWrEn ? sbWrMask : T_828;
  assign T_830 = dbRamWrEn | dbRamRdEn;
  assign T_831 = sbRamRdEn | sbRamWrEn;
  assign T_832 = T_830 & T_831;
  assign T_834 = T_832 == 1'h0;
  assign T_835 = T_834 | reset;
  assign T_837 = T_835 == 1'h0;
  assign dbRamWrDataVec = {dbRamWrData,dbRamWrData};
  assign T_838 = ramWrMask & sbRamWrData;
  assign T_839 = ~ ramWrMask;
  assign T_840 = T_839 & ramRdData;
  assign T_841 = T_838 | T_840;
  assign T_842 = ramWrMask & dbRamWrDataVec;
  assign T_845 = T_842 | T_840;
  assign T_846 = sbRamWrEn ? T_841 : T_845;
  assign T_847 = sbRamWrEn | sbRamRdEn;
  assign T_848 = dbRamAddr[2:1];
  assign T_849 = T_847 ? sbRamAddr : T_848;
  assign T_852 = sbRamWrEn | dbRamWrEn;
  assign T_875_interrupt = T_895;
  assign T_875_haltnot = T_894;
  assign T_875_reserved0 = T_893;
  assign T_875_buserror = T_892;
  assign T_875_serial = T_891;
  assign T_875_autoincrement = T_890;
  assign T_875_access = T_889;
  assign T_875_hartid = T_888;
  assign T_875_ndreset = T_887;
  assign T_875_fullreset = T_886;
  assign T_886 = dbReq_data[0];
  assign T_887 = dbReq_data[1];
  assign T_888 = dbReq_data[11:2];
  assign T_889 = dbReq_data[14:12];
  assign T_890 = dbReq_data[15];
  assign T_891 = dbReq_data[18:16];
  assign T_892 = dbReq_data[21:19];
  assign T_893 = dbReq_data[31:22];
  assign T_894 = dbReq_data[32];
  assign T_895 = dbReq_data[33];
  assign T_904_interrupt = T_895;
  assign T_904_haltnot = T_894;
  assign T_904_data = T_908;
  assign T_908 = dbReq_data[31:0];
  assign T_913 = dbReq_addr[4:4];
  assign T_915 = T_913 == 1'h0;
  assign GEN_31 = T_915 ? dbWrEn : 1'h0;
  assign T_917 = dbReq_addr == 5'h10;
  assign T_919 = T_915 == 1'h0;
  assign T_920 = T_919 & T_917;
  assign GEN_32 = T_920 ? dbWrEn : 1'h0;
  assign T_924 = T_917 == 1'h0;
  assign T_925 = T_919 & T_924;
  assign GEN_33 = reset ? CONTROLReset_interrupt : CONTROLReg_interrupt;
  assign GEN_34 = reset ? CONTROLReset_haltnot : CONTROLReg_haltnot;
  assign GEN_35 = reset ? CONTROLReset_reserved0 : CONTROLReg_reserved0;
  assign GEN_36 = reset ? CONTROLReset_buserror : CONTROLReg_buserror;
  assign GEN_37 = reset ? CONTROLReset_serial : CONTROLReg_serial;
  assign GEN_38 = reset ? CONTROLReset_autoincrement : CONTROLReg_autoincrement;
  assign GEN_39 = reset ? CONTROLReset_access : CONTROLReg_access;
  assign GEN_40 = reset ? CONTROLReset_hartid : CONTROLReg_hartid;
  assign GEN_41 = reset ? CONTROLReset_ndreset : CONTROLReg_ndreset;
  assign GEN_42 = reset ? CONTROLReset_fullreset : CONTROLReg_fullreset;
  assign GEN_43 = reset ? 1'h0 : ndresetCtrReg;
  assign T_928 = reset == 1'h0;
  assign T_929 = T_928 & CONTROLWrEn;
  assign T_930 = CONTROLReg_fullreset | CONTROLWrData_fullreset;
  assign GEN_44 = CONTROLWrData_ndreset ? 1'h1 : GEN_43;
  assign T_933 = CONTROLWrData_ndreset == 1'h0;
  assign T_935 = ndresetCtrReg == 1'h0;
  assign T_938 = ndresetCtrReg - 1'h1;
  assign T_939 = T_938[0:0];
  assign T_940 = T_935 ? 1'h0 : T_939;
  assign GEN_45 = T_933 ? T_940 : GEN_44;
  assign GEN_46 = T_929 ? CONTROLWrData_hartid : GEN_40;
  assign GEN_47 = T_929 ? T_930 : GEN_42;
  assign GEN_48 = T_929 ? GEN_45 : GEN_43;
  assign T_945 = T_928 & T_723;
  assign GEN_49 = T_945 ? T_940 : GEN_48;
  assign GEN_2 = interruptRegs_0;
  assign GEN_3 = haltnotRegs_0;
  assign GEN_4 = interruptRegs_0;
  assign GEN_5 = haltnotRegs_0;
  assign T_958 = dbReq_addr == 5'h0;
  assign GEN_50 = T_958 ? haltnotStatus_0 : 32'h0;
  assign T_963 = {RAMRdData_interrupt,RAMRdData_haltnot};
  assign T_964 = {T_963,RAMRdData_data};
  assign GEN_51 = T_915 ? T_964 : 34'h0;
  assign T_970 = {CONTROLRdData_ndreset,CONTROLRdData_fullreset};
  assign T_971 = {CONTROLRdData_autoincrement,CONTROLRdData_access};
  assign T_972 = {T_971,CONTROLRdData_hartid};
  assign T_973 = {T_972,T_970};
  assign T_974 = {CONTROLRdData_buserror,CONTROLRdData_serial};
  assign T_975 = {CONTROLRdData_interrupt,CONTROLRdData_haltnot};
  assign T_976 = {T_975,CONTROLRdData_reserved0};
  assign T_977 = {T_976,T_974};
  assign T_978 = {T_977,T_973};
  assign GEN_53 = T_920 ? T_978 : GEN_51;
  assign T_980 = dbReq_addr == 5'h11;
  assign T_986 = T_925 & T_980;
  assign T_987 = {DMINFORdData_authbusy,DMINFORdData_authtype};
  assign T_988 = {T_987,DMINFORdData_version};
  assign T_989 = {DMINFORdData_reserved1,DMINFORdData_authenticated};
  assign T_990 = {DMINFORdData_dramsize,DMINFORdData_haltsum};
  assign T_991 = {T_990,T_989};
  assign T_992 = {T_991,T_988};
  assign T_993 = {DMINFORdData_access16,DMINFORdData_accesss8};
  assign T_994 = {DMINFORdData_access64,DMINFORdData_access32};
  assign T_995 = {T_994,T_993};
  assign T_996 = {DMINFORdData_serialcount,DMINFORdData_access128};
  assign T_997 = {DMINFORdData_reserved0,DMINFORdData_abussize};
  assign T_998 = {T_997,T_996};
  assign T_999 = {T_998,T_995};
  assign T_1000 = {T_999,T_992};
  assign GEN_54 = T_986 ? T_1000 : GEN_53;
  assign T_1002 = dbReq_addr == 5'h1b;
  assign T_1009 = T_980 == 1'h0;
  assign T_1010 = T_925 & T_1009;
  assign T_1011 = T_1010 & T_1002;
  assign GEN_55 = T_1011 ? 34'h0 : GEN_54;
  assign T_1013 = dbReq_addr[4:2];
  assign T_1015 = T_1013 == 3'h7;
  assign T_1025 = T_1002 == 1'h0;
  assign T_1026 = T_1010 & T_1025;
  assign T_1027 = T_1026 & T_1015;
  assign GEN_56 = T_1027 ? {{2'd0}, rdHaltnotStatus} : GEN_55;
  assign T_1040 = T_1015 == 1'h0;
  assign T_1041 = T_1026 & T_1040;
  assign GEN_57 = T_1041 ? 34'h0 : GEN_56;
  assign T_1043 = dbRdData[33];
  assign T_1045 = dbReq_op == 2'h3;
  assign T_1046 = T_1043 & T_1045;
  assign T_1048 = dbReq_op == 2'h2;
  assign T_1051 = ~ rdCondWrFailure;
  assign T_1052 = T_1045 & T_1051;
  assign T_1053 = T_1048 | T_1052;
  assign T_1056 = rdCondWrFailure ? 2'h1 : 2'h0;
  assign T_1058 = stallFromSb == 1'h0;
  assign T_1059 = dbStateReg == 1'h0;
  assign T_1061 = io_db_resp_ready & io_db_resp_valid;
  assign T_1062 = dbStateReg & T_1061;
  assign T_1063 = T_1059 | T_1062;
  assign T_1064 = T_1058 & T_1063;
  assign T_1066 = io_db_req_ready & io_db_req_valid;
  assign T_1068 = dbWrNeeded & T_1066;
  assign GEN_58 = T_1066 ? 1'h1 : dbStateReg;
  assign GEN_59 = T_1066 ? dbResult_resp : dbRespReg_resp;
  assign GEN_60 = T_1066 ? dbResult_data : dbRespReg_data;
  assign GEN_61 = T_1059 ? GEN_58 : dbStateReg;
  assign GEN_62 = T_1059 ? GEN_59 : dbRespReg_resp;
  assign GEN_63 = T_1059 ? GEN_60 : dbRespReg_data;
  assign T_1073 = T_1059 == 1'h0;
  assign T_1074 = T_1073 & dbStateReg;
  assign GEN_64 = T_1066 ? 1'h1 : GEN_61;
  assign GEN_65 = T_1066 ? dbResult_resp : GEN_62;
  assign GEN_66 = T_1066 ? dbResult_data : GEN_63;
  assign T_1078 = T_1066 == 1'h0;
  assign T_1079 = T_1078 & T_1061;
  assign GEN_67 = T_1079 ? 1'h0 : GEN_64;
  assign GEN_68 = T_1074 ? GEN_67 : GEN_61;
  assign GEN_69 = T_1074 ? GEN_65 : GEN_62;
  assign GEN_70 = T_1074 ? GEN_66 : GEN_63;
  assign T_1101_0 = 64'hc0006f03c0006f;
  assign T_1101_1 = 64'h80006ffff00413;
  assign T_1101_2 = 64'hff0000f00000413;
  assign T_1101_3 = 64'h40802c2341802483;
  assign T_1101_4 = 64'h10802023f1402473;
  assign T_1101_5 = 64'h8474137b002473;
  assign T_1101_6 = 64'h7b20247302041a63;
  assign T_1101_7 = 64'h7b2410737b200073;
  assign T_1101_8 = 64'h1c0474137b002473;
  assign T_1101_9 = 64'h41663f4040413;
  assign T_1101_10 = 64'h4000006740902c23;
  assign T_1101_11 = 64'h10802623f1402473;
  assign T_1101_12 = 64'h7b0024737b046073;
  assign T_1101_13 = 64'hfe040ce302047413;
  assign T_1101_14 = 64'hfe1ff06f;
  assign T_1104 = T_1105;
  assign T_1105 = sbAddr[6:3];
  assign GEN_6 = GEN_84;
  assign GEN_71 = 4'h1 == T_1104 ? T_1101_1 : T_1101_0;
  assign GEN_72 = 4'h2 == T_1104 ? T_1101_2 : GEN_71;
  assign GEN_73 = 4'h3 == T_1104 ? T_1101_3 : GEN_72;
  assign GEN_74 = 4'h4 == T_1104 ? T_1101_4 : GEN_73;
  assign GEN_75 = 4'h5 == T_1104 ? T_1101_5 : GEN_74;
  assign GEN_76 = 4'h6 == T_1104 ? T_1101_6 : GEN_75;
  assign GEN_77 = 4'h7 == T_1104 ? T_1101_7 : GEN_76;
  assign GEN_78 = 4'h8 == T_1104 ? T_1101_8 : GEN_77;
  assign GEN_79 = 4'h9 == T_1104 ? T_1101_9 : GEN_78;
  assign GEN_80 = 4'ha == T_1104 ? T_1101_10 : GEN_79;
  assign GEN_81 = 4'hb == T_1104 ? T_1101_11 : GEN_80;
  assign GEN_82 = 4'hc == T_1104 ? T_1101_12 : GEN_81;
  assign GEN_83 = 4'hd == T_1104 ? T_1101_13 : GEN_82;
  assign GEN_84 = 4'he == T_1104 ? T_1101_14 : GEN_83;
  assign T_1109 = sbWrData[31:0];
  assign T_1110 = sbWrData[63:32];
  assign T_1116_0 = T_1109;
  assign T_1116_1 = T_1110;
  assign T_1118 = sbWrMask[31:0];
  assign T_1119 = sbWrMask[63:32];
  assign T_1125_0 = T_1118;
  assign T_1125_1 = T_1119;
  assign GEN_7 = T_1116_1;
  assign GEN_8 = T_1116_0;
  assign T_1131 = sbAddr[11:8];
  assign T_1133 = T_1131 == 4'h4;
  assign GEN_87 = T_1133 ? sbWrEn : 1'h0;
  assign T_1134 = sbAddr[11:3];
  assign T_1137 = T_1134 == 9'h21;
  assign GEN_9 = T_1125_1;
  assign T_1141 = GEN_9 != 32'h0;
  assign T_1142 = T_1137 & T_1141;
  assign T_1143 = T_1142 & sbWrEn;
  assign T_1147 = T_1134 == 9'h20;
  assign GEN_10 = T_1125_0;
  assign T_1151 = GEN_10 != 32'h0;
  assign T_1152 = T_1147 & T_1151;
  assign T_1153 = T_1152 & sbWrEn;
  assign GEN_91 = T_1133 ? sbRamRdData : 64'h0;
  assign GEN_92 = T_1133 ? sbRdEn : 1'h0;
  assign T_1162 = T_1131 == 4'h8;
  assign T_1165 = T_1131 == 4'h9;
  assign T_1166 = T_1162 | T_1165;
  assign T_1168 = T_1133 == 1'h0;
  assign T_1169 = T_1168 & T_1166;
  assign GEN_93 = T_1169 ? sbRomRdData : GEN_91;
  assign T_1173 = T_1166 == 1'h0;
  assign T_1174 = T_1168 & T_1173;
  assign GEN_94 = T_1174 ? 64'h0 : GEN_93;
  assign T_1203 = sbAcqReg_a_type == 3'h0;
  assign sbReg_get = sbAcqReg_is_builtin_type & T_1203;
  assign T_1204 = sbAcqReg_a_type == 3'h1;
  assign sbReg_getblk = sbAcqReg_is_builtin_type & T_1204;
  assign T_1205 = sbAcqReg_a_type == 3'h2;
  assign sbReg_put = sbAcqReg_is_builtin_type & T_1205;
  assign T_1206 = sbAcqReg_a_type == 3'h3;
  assign sbReg_putblk = sbAcqReg_is_builtin_type & T_1206;
  assign sbMultibeat = sbReg_getblk & sbAcqValidReg;
  assign T_1208 = sbAcqReg_addr_beat + 3'h1;
  assign sbBeatInc1 = T_1208[2:0];
  assign sbLast = sbAcqReg_addr_beat == 3'h7;
  assign T_1217_0 = 3'h0;
  assign T_1217_1 = 3'h4;
  assign T_1219 = sbAcqReg_a_type == T_1217_0;
  assign T_1220 = sbAcqReg_a_type == T_1217_1;
  assign T_1221 = T_1219 | T_1220;
  assign T_1222 = sbAcqReg_is_builtin_type & T_1221;
  assign T_1223 = sbAcqReg_union[11:9];
  assign T_1225 = T_1222 ? T_1223 : 3'h0;
  assign T_1226 = {sbAcqReg_addr_block,sbAcqReg_addr_beat};
  assign T_1227 = {T_1226,T_1225};
  assign T_1228 = sbReg_get | sbReg_getblk;
  assign T_1229 = sbAcqValidReg & T_1228;
  assign T_1230 = sbReg_put | sbReg_putblk;
  assign T_1231 = sbAcqValidReg & T_1230;
  assign T_1233 = sbAcqReg_a_type == 3'h4;
  assign T_1234 = sbAcqReg_is_builtin_type & T_1233;
  assign T_1236 = T_1223[2];
  assign T_1238 = 2'h1 << T_1236;
  assign T_1239 = T_1238[0];
  assign T_1240 = T_1238[1];
  assign T_1244 = T_1239 ? 4'hf : 4'h0;
  assign T_1248 = T_1240 ? 4'hf : 4'h0;
  assign T_1249 = {T_1248,T_1244};
  assign T_1256 = sbReg_putblk | sbReg_put;
  assign T_1257 = sbAcqReg_union[8:1];
  assign T_1259 = T_1256 ? T_1257 : 8'h0;
  assign T_1260 = T_1234 ? T_1249 : T_1259;
  assign T_1261 = T_1260[0];
  assign T_1262 = T_1260[1];
  assign T_1263 = T_1260[2];
  assign T_1264 = T_1260[3];
  assign T_1265 = T_1260[4];
  assign T_1266 = T_1260[5];
  assign T_1267 = T_1260[6];
  assign T_1268 = T_1260[7];
  assign T_1272 = T_1261 ? 8'hff : 8'h0;
  assign T_1276 = T_1262 ? 8'hff : 8'h0;
  assign T_1280 = T_1263 ? 8'hff : 8'h0;
  assign T_1284 = T_1264 ? 8'hff : 8'h0;
  assign T_1288 = T_1265 ? 8'hff : 8'h0;
  assign T_1292 = T_1266 ? 8'hff : 8'h0;
  assign T_1296 = T_1267 ? 8'hff : 8'h0;
  assign T_1300 = T_1268 ? 8'hff : 8'h0;
  assign T_1301 = {T_1276,T_1272};
  assign T_1302 = {T_1284,T_1280};
  assign T_1303 = {T_1302,T_1301};
  assign T_1304 = {T_1292,T_1288};
  assign T_1305 = {T_1300,T_1296};
  assign T_1306 = {T_1305,T_1304};
  assign T_1307 = {T_1306,T_1303};
  assign T_1308 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign GEN_95 = T_1308 ? io_tl_acquire_bits_addr_block : sbAcqReg_addr_block;
  assign GEN_96 = T_1308 ? io_tl_acquire_bits_client_xact_id : sbAcqReg_client_xact_id;
  assign GEN_97 = T_1308 ? io_tl_acquire_bits_addr_beat : sbAcqReg_addr_beat;
  assign GEN_98 = T_1308 ? io_tl_acquire_bits_is_builtin_type : sbAcqReg_is_builtin_type;
  assign GEN_99 = T_1308 ? io_tl_acquire_bits_a_type : sbAcqReg_a_type;
  assign GEN_100 = T_1308 ? io_tl_acquire_bits_union : sbAcqReg_union;
  assign GEN_101 = T_1308 ? io_tl_acquire_bits_data : sbAcqReg_data;
  assign GEN_102 = T_1308 ? 1'h1 : sbAcqValidReg;
  assign T_1310 = io_tl_grant_ready & io_tl_grant_valid;
  assign T_1312 = T_1308 == 1'h0;
  assign T_1313 = T_1312 & T_1310;
  assign GEN_103 = sbLast ? 1'h0 : GEN_102;
  assign GEN_104 = sbMultibeat ? sbBeatInc1 : GEN_97;
  assign GEN_105 = sbMultibeat ? GEN_103 : GEN_102;
  assign T_1316 = sbMultibeat == 1'h0;
  assign GEN_106 = T_1316 ? 1'h0 : GEN_105;
  assign GEN_107 = T_1313 ? GEN_104 : GEN_97;
  assign GEN_108 = T_1313 ? GEN_106 : GEN_102;
  assign T_1334 = 3'h6 == sbAcqReg_a_type;
  assign T_1335 = T_1334 ? 3'h1 : 3'h3;
  assign T_1336 = 3'h5 == sbAcqReg_a_type;
  assign T_1337 = T_1336 ? 3'h1 : T_1335;
  assign T_1338 = 3'h4 == sbAcqReg_a_type;
  assign T_1339 = T_1338 ? 3'h4 : T_1337;
  assign T_1340 = 3'h3 == sbAcqReg_a_type;
  assign T_1341 = T_1340 ? 3'h3 : T_1339;
  assign T_1342 = 3'h2 == sbAcqReg_a_type;
  assign T_1343 = T_1342 ? 3'h3 : T_1341;
  assign T_1344 = 3'h1 == sbAcqReg_a_type;
  assign T_1345 = T_1344 ? 3'h5 : T_1343;
  assign T_1346 = 3'h0 == sbAcqReg_a_type;
  assign T_1347 = T_1346 ? 3'h4 : T_1345;
  assign T_1371_addr_beat = sbAcqReg_addr_beat;
  assign T_1371_client_xact_id = sbAcqReg_client_xact_id;
  assign T_1371_manager_xact_id = 1'h0;
  assign T_1371_is_builtin_type = 1'h1;
  assign T_1371_g_type = {{1'd0}, T_1347};
  assign T_1371_data = sbRdData;
  assign T_1396 = sbLast == 1'h0;
  assign T_1397 = sbMultibeat & T_1396;
  assign T_1399 = io_tl_grant_ready == 1'h0;
  assign T_1400 = io_tl_grant_valid & T_1399;
  assign T_1401 = T_1397 | T_1400;
  assign sbStall = T_1401 | stallFromDb;
  assign T_1403 = sbStall == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_26 = {1{$random}};
  CONTROLReg_interrupt = GEN_26[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_27 = {1{$random}};
  CONTROLReg_haltnot = GEN_27[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_28 = {1{$random}};
  CONTROLReg_reserved0 = GEN_28[9:0];
  `endif
  `ifdef RANDOMIZE
  GEN_29 = {1{$random}};
  CONTROLReg_buserror = GEN_29[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_30 = {1{$random}};
  CONTROLReg_serial = GEN_30[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_52 = {1{$random}};
  CONTROLReg_autoincrement = GEN_52[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_85 = {1{$random}};
  CONTROLReg_access = GEN_85[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_86 = {1{$random}};
  CONTROLReg_hartid = GEN_86[9:0];
  `endif
  `ifdef RANDOMIZE
  GEN_88 = {1{$random}};
  CONTROLReg_ndreset = GEN_88[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_89 = {1{$random}};
  CONTROLReg_fullreset = GEN_89[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_90 = {1{$random}};
  ndresetCtrReg = GEN_90[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_109 = {1{$random}};
  interruptRegs_0 = GEN_109[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_110 = {1{$random}};
  haltnotRegs_0 = GEN_110[0:0];
  `endif
  GEN_111 = {2{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ramMem[initvar] = GEN_111[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_112 = {1{$random}};
  dbStateReg = GEN_112[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_113 = {1{$random}};
  dbRespReg_resp = GEN_113[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_114 = {2{$random}};
  dbRespReg_data = GEN_114[33:0];
  `endif
  `ifdef RANDOMIZE
  GEN_115 = {1{$random}};
  sbAcqReg_addr_block = GEN_115[25:0];
  `endif
  `ifdef RANDOMIZE
  GEN_116 = {1{$random}};
  sbAcqReg_client_xact_id = GEN_116[1:0];
  `endif
  `ifdef RANDOMIZE
  GEN_117 = {1{$random}};
  sbAcqReg_addr_beat = GEN_117[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_118 = {1{$random}};
  sbAcqReg_is_builtin_type = GEN_118[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_119 = {1{$random}};
  sbAcqReg_a_type = GEN_119[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_120 = {1{$random}};
  sbAcqReg_union = GEN_120[11:0];
  `endif
  `ifdef RANDOMIZE
  GEN_121 = {2{$random}};
  sbAcqReg_data = GEN_121[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_122 = {1{$random}};
  sbAcqValidReg = GEN_122[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_interrupt <= CONTROLReset_interrupt;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_haltnot <= CONTROLReset_haltnot;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_reserved0 <= CONTROLReset_reserved0;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_buserror <= CONTROLReset_buserror;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_serial <= CONTROLReset_serial;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_autoincrement <= CONTROLReset_autoincrement;
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_access <= CONTROLReset_access;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_929) begin
        CONTROLReg_hartid <= CONTROLWrData_hartid;
      end else begin
        if(reset) begin
          CONTROLReg_hartid <= CONTROLReset_hartid;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(reset) begin
        CONTROLReg_ndreset <= CONTROLReset_ndreset;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_929) begin
        CONTROLReg_fullreset <= T_930;
      end else begin
        if(reset) begin
          CONTROLReg_fullreset <= CONTROLReset_fullreset;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_945) begin
        if(T_935) begin
          ndresetCtrReg <= 1'h0;
        end else begin
          ndresetCtrReg <= T_939;
        end
      end else begin
        if(T_929) begin
          if(T_933) begin
            if(T_935) begin
              ndresetCtrReg <= 1'h0;
            end else begin
              ndresetCtrReg <= T_939;
            end
          end else begin
            if(CONTROLWrData_ndreset) begin
              ndresetCtrReg <= 1'h1;
            end else begin
              if(reset) begin
                ndresetCtrReg <= 1'h0;
              end
            end
          end
        end else begin
          if(reset) begin
            ndresetCtrReg <= 1'h0;
          end
        end
      end
    end
    if(reset) begin
      interruptRegs_0 <= T_655_0;
    end else begin
      if(T_733) begin
        if(T_735) begin
          interruptRegs_0 <= 1'h0;
        end else begin
          if(T_724) begin
            if(T_726) begin
              interruptRegs_0 <= T_727;
            end else begin
              if(CONTROLWrEn) begin
                if(T_720) begin
                  interruptRegs_0 <= T_721;
                end
              end
            end
          end else begin
            if(CONTROLWrEn) begin
              if(T_720) begin
                interruptRegs_0 <= T_721;
              end
            end
          end
        end
      end else begin
        if(T_724) begin
          if(T_726) begin
            interruptRegs_0 <= T_727;
          end else begin
            if(CONTROLWrEn) begin
              if(T_720) begin
                interruptRegs_0 <= T_721;
              end
            end
          end
        end else begin
          if(CONTROLWrEn) begin
            if(T_720) begin
              interruptRegs_0 <= T_721;
            end
          end
        end
      end
    end
    if(reset) begin
      haltnotRegs_0 <= T_666_0;
    end else begin
      if(T_751) begin
        if(T_726) begin
          haltnotRegs_0 <= T_754;
        end else begin
          if(T_742) begin
            if(T_720) begin
              haltnotRegs_0 <= T_745;
            end else begin
              if(SETHALTNOTWrEn) begin
                if(T_738) begin
                  haltnotRegs_0 <= 1'h1;
                end
              end
            end
          end else begin
            if(SETHALTNOTWrEn) begin
              if(T_738) begin
                haltnotRegs_0 <= 1'h1;
              end
            end
          end
        end
      end else begin
        if(T_742) begin
          if(T_720) begin
            haltnotRegs_0 <= T_745;
          end else begin
            if(SETHALTNOTWrEn) begin
              if(T_738) begin
                haltnotRegs_0 <= 1'h1;
              end
            end
          end
        end else begin
          if(SETHALTNOTWrEn) begin
            if(T_738) begin
              haltnotRegs_0 <= 1'h1;
            end
          end
        end
      end
    end
    if(ramMem_T_851_en & ramMem_T_851_mask) begin
      ramMem[ramMem_T_851_addr] <= ramMem_T_851_data;
    end
    if(reset) begin
      dbStateReg <= 1'h0;
    end else begin
      if(T_1074) begin
        if(T_1079) begin
          dbStateReg <= 1'h0;
        end else begin
          if(T_1066) begin
            dbStateReg <= 1'h1;
          end else begin
            if(T_1059) begin
              if(T_1066) begin
                dbStateReg <= 1'h1;
              end
            end
          end
        end
      end else begin
        if(T_1059) begin
          if(T_1066) begin
            dbStateReg <= 1'h1;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1074) begin
        if(T_1066) begin
          dbRespReg_resp <= dbResult_resp;
        end else begin
          if(T_1059) begin
            if(T_1066) begin
              dbRespReg_resp <= dbResult_resp;
            end
          end
        end
      end else begin
        if(T_1059) begin
          if(T_1066) begin
            dbRespReg_resp <= dbResult_resp;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1074) begin
        if(T_1066) begin
          dbRespReg_data <= dbResult_data;
        end else begin
          if(T_1059) begin
            if(T_1066) begin
              dbRespReg_data <= dbResult_data;
            end
          end
        end
      end else begin
        if(T_1059) begin
          if(T_1066) begin
            dbRespReg_data <= dbResult_data;
          end
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1308) begin
        sbAcqReg_addr_block <= io_tl_acquire_bits_addr_block;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1308) begin
        sbAcqReg_client_xact_id <= io_tl_acquire_bits_client_xact_id;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1313) begin
        if(sbMultibeat) begin
          sbAcqReg_addr_beat <= sbBeatInc1;
        end else begin
          if(T_1308) begin
            sbAcqReg_addr_beat <= io_tl_acquire_bits_addr_beat;
          end
        end
      end else begin
        if(T_1308) begin
          sbAcqReg_addr_beat <= io_tl_acquire_bits_addr_beat;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1308) begin
        sbAcqReg_is_builtin_type <= io_tl_acquire_bits_is_builtin_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1308) begin
        sbAcqReg_a_type <= io_tl_acquire_bits_a_type;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1308) begin
        sbAcqReg_union <= io_tl_acquire_bits_union;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1308) begin
        sbAcqReg_data <= io_tl_acquire_bits_data;
      end
    end
    if(reset) begin
      sbAcqValidReg <= 1'h0;
    end else begin
      if(T_1313) begin
        if(T_1316) begin
          sbAcqValidReg <= 1'h0;
        end else begin
          if(sbMultibeat) begin
            if(sbLast) begin
              sbAcqValidReg <= 1'h0;
            end else begin
              if(T_1308) begin
                sbAcqValidReg <= 1'h1;
              end
            end
          end else begin
            if(T_1308) begin
              sbAcqValidReg <= 1'h1;
            end
          end
        end
      end else begin
        if(T_1308) begin
          sbAcqValidReg <= 1'h1;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_837) begin
          $fwrite(32'h80000002,"Assertion failed: Stall logic should have prevented concurrent SB/DB RAM Access\n    at Debug.scala:652 assert (!((dbRamWrEn | dbRamRdEn) & (sbRamRdEn | sbRamWrEn)), ---Stall logic should have prevented concurrent SB/DB RAM Access---)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_837) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module PRCI(
  input   clk,
  input   reset,
  input   io_interrupts_0_meip,
  input   io_interrupts_0_seip,
  input   io_interrupts_0_debug,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [11:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data,
  output  io_tiles_0_reset,
  output  io_tiles_0_id,
  output  io_tiles_0_interrupts_meip,
  output  io_tiles_0_interrupts_seip,
  output  io_tiles_0_interrupts_debug,
  output  io_tiles_0_interrupts_mtip,
  output  io_tiles_0_interrupts_msip,
  input   io_rtcTick
);
  reg [63:0] timecmp_0;
  reg [63:0] GEN_2;
  reg [63:0] time$;
  reg [63:0] GEN_3;
  wire [64:0] T_525;
  wire [63:0] T_526;
  wire [63:0] GEN_0;
  wire [31:0] T_533_0;
  reg [31:0] ipi_0;
  reg [31:0] GEN_6;
  wire  acq_clk;
  wire  acq_reset;
  wire  acq_io_enq_ready;
  wire  acq_io_enq_valid;
  wire [25:0] acq_io_enq_bits_addr_block;
  wire [1:0] acq_io_enq_bits_client_xact_id;
  wire [2:0] acq_io_enq_bits_addr_beat;
  wire  acq_io_enq_bits_is_builtin_type;
  wire [2:0] acq_io_enq_bits_a_type;
  wire [11:0] acq_io_enq_bits_union;
  wire [63:0] acq_io_enq_bits_data;
  wire  acq_io_deq_ready;
  wire  acq_io_deq_valid;
  wire [25:0] acq_io_deq_bits_addr_block;
  wire [1:0] acq_io_deq_bits_client_xact_id;
  wire [2:0] acq_io_deq_bits_addr_beat;
  wire  acq_io_deq_bits_is_builtin_type;
  wire [2:0] acq_io_deq_bits_a_type;
  wire [11:0] acq_io_deq_bits_union;
  wire [63:0] acq_io_deq_bits_data;
  wire  acq_io_count;
  wire [2:0] T_568_0;
  wire [2:0] T_568_1;
  wire  T_570;
  wire  T_571;
  wire  T_572;
  wire  T_573;
  wire [2:0] T_574;
  wire [2:0] T_576;
  wire [28:0] T_577;
  wire [31:0] T_578;
  wire [15:0] addr;
  wire [63:0] rdata;
  wire  T_598;
  wire [2:0] T_599;
  wire  T_600;
  wire [2:0] T_601;
  wire  T_602;
  wire [2:0] T_603;
  wire  T_604;
  wire [2:0] T_605;
  wire  T_606;
  wire [2:0] T_607;
  wire  T_608;
  wire [2:0] T_609;
  wire  T_610;
  wire [2:0] T_611;
  wire [2:0] T_636_addr_beat;
  wire [1:0] T_636_client_xact_id;
  wire  T_636_manager_xact_id;
  wire  T_636_is_builtin_type;
  wire [3:0] T_636_g_type;
  wire [63:0] T_636_data;
  wire  T_658;
  wire [64:0] T_660;
  wire [63:0] T_661;
  wire [63:0] T_667_0;
  wire [2:0] T_676_0;
  wire [2:0] T_676_1;
  wire [63:0] GEN_4;
  wire  T_688;
  wire  T_690;
  wire  T_691;
  wire [2:0] T_699_0;
  wire [2:0] T_699_1;
  wire [2:0] T_717_0;
  wire [2:0] T_717_1;
  wire  T_729;
  wire  T_730;
  wire  T_732;
  wire [1:0] T_734;
  wire  T_735;
  wire  T_736;
  wire [3:0] T_740;
  wire [3:0] T_744;
  wire [7:0] T_745;
  wire  T_747;
  wire  T_748;
  wire  T_750;
  wire  T_751;
  wire  T_752;
  wire [7:0] T_753;
  wire [7:0] T_755;
  wire [7:0] T_756;
  wire  T_757;
  wire  T_758;
  wire  T_759;
  wire  T_760;
  wire  T_761;
  wire  T_762;
  wire  T_763;
  wire  T_764;
  wire [7:0] T_768;
  wire [7:0] T_772;
  wire [7:0] T_776;
  wire [7:0] T_780;
  wire [7:0] T_784;
  wire [7:0] T_788;
  wire [7:0] T_792;
  wire [7:0] T_796;
  wire [15:0] T_797;
  wire [15:0] T_798;
  wire [31:0] T_799;
  wire [15:0] T_800;
  wire [15:0] T_801;
  wire [31:0] T_802;
  wire [63:0] T_803;
  wire [63:0] T_804;
  wire [63:0] T_881;
  wire [63:0] T_882;
  wire [63:0] T_883;
  wire [63:0] GEN_5;
  wire [63:0] GEN_10;
  wire [63:0] GEN_11;
  wire  T_895;
  wire  T_896;
  wire [2:0] T_904_0;
  wire [2:0] T_904_1;
  wire [2:0] T_922_0;
  wire [2:0] T_922_1;
  wire [63:0] GEN_19;
  wire [63:0] T_1087;
  wire [63:0] T_1088;
  wire [63:0] GEN_12;
  wire [63:0] T_1099;
  wire [63:0] GEN_17;
  wire [63:0] GEN_18;
  wire  T_1100;
  wire  T_1101;
  reg  GEN_1;
  reg [31:0] GEN_7;
  Queue_8 acq (
    .clk(acq_clk),
    .reset(acq_reset),
    .io_enq_ready(acq_io_enq_ready),
    .io_enq_valid(acq_io_enq_valid),
    .io_enq_bits_addr_block(acq_io_enq_bits_addr_block),
    .io_enq_bits_client_xact_id(acq_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(acq_io_enq_bits_addr_beat),
    .io_enq_bits_is_builtin_type(acq_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(acq_io_enq_bits_a_type),
    .io_enq_bits_union(acq_io_enq_bits_union),
    .io_enq_bits_data(acq_io_enq_bits_data),
    .io_deq_ready(acq_io_deq_ready),
    .io_deq_valid(acq_io_deq_valid),
    .io_deq_bits_addr_block(acq_io_deq_bits_addr_block),
    .io_deq_bits_client_xact_id(acq_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(acq_io_deq_bits_addr_beat),
    .io_deq_bits_is_builtin_type(acq_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(acq_io_deq_bits_a_type),
    .io_deq_bits_union(acq_io_deq_bits_union),
    .io_deq_bits_data(acq_io_deq_bits_data),
    .io_count(acq_io_count)
  );
  assign io_tl_acquire_ready = acq_io_enq_ready;
  assign io_tl_grant_valid = acq_io_deq_valid;
  assign io_tl_grant_bits_addr_beat = T_636_addr_beat;
  assign io_tl_grant_bits_client_xact_id = T_636_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = T_636_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = T_636_is_builtin_type;
  assign io_tl_grant_bits_g_type = T_636_g_type;
  assign io_tl_grant_bits_data = T_636_data;
  assign io_tiles_0_reset = GEN_1;
  assign io_tiles_0_id = 1'h0;
  assign io_tiles_0_interrupts_meip = io_interrupts_0_meip;
  assign io_tiles_0_interrupts_seip = io_interrupts_0_seip;
  assign io_tiles_0_interrupts_debug = io_interrupts_0_debug;
  assign io_tiles_0_interrupts_mtip = T_1101;
  assign io_tiles_0_interrupts_msip = T_1100;
  assign T_525 = time$ + 64'h1;
  assign T_526 = T_525[63:0];
  assign GEN_0 = io_rtcTick ? T_526 : time$;
  assign T_533_0 = 32'h0;
  assign acq_clk = clk;
  assign acq_reset = reset;
  assign acq_io_enq_valid = io_tl_acquire_valid;
  assign acq_io_enq_bits_addr_block = io_tl_acquire_bits_addr_block;
  assign acq_io_enq_bits_client_xact_id = io_tl_acquire_bits_client_xact_id;
  assign acq_io_enq_bits_addr_beat = io_tl_acquire_bits_addr_beat;
  assign acq_io_enq_bits_is_builtin_type = io_tl_acquire_bits_is_builtin_type;
  assign acq_io_enq_bits_a_type = io_tl_acquire_bits_a_type;
  assign acq_io_enq_bits_union = io_tl_acquire_bits_union;
  assign acq_io_enq_bits_data = io_tl_acquire_bits_data;
  assign acq_io_deq_ready = io_tl_grant_ready;
  assign T_568_0 = 3'h0;
  assign T_568_1 = 3'h4;
  assign T_570 = acq_io_deq_bits_a_type == T_568_0;
  assign T_571 = acq_io_deq_bits_a_type == T_568_1;
  assign T_572 = T_570 | T_571;
  assign T_573 = acq_io_deq_bits_is_builtin_type & T_572;
  assign T_574 = acq_io_deq_bits_union[11:9];
  assign T_576 = T_573 ? T_574 : 3'h0;
  assign T_577 = {acq_io_deq_bits_addr_block,acq_io_deq_bits_addr_beat};
  assign T_578 = {T_577,T_576};
  assign addr = T_578[15:0];
  assign rdata = GEN_18;
  assign T_598 = 3'h6 == acq_io_deq_bits_a_type;
  assign T_599 = T_598 ? 3'h1 : 3'h3;
  assign T_600 = 3'h5 == acq_io_deq_bits_a_type;
  assign T_601 = T_600 ? 3'h1 : T_599;
  assign T_602 = 3'h4 == acq_io_deq_bits_a_type;
  assign T_603 = T_602 ? 3'h4 : T_601;
  assign T_604 = 3'h3 == acq_io_deq_bits_a_type;
  assign T_605 = T_604 ? 3'h3 : T_603;
  assign T_606 = 3'h2 == acq_io_deq_bits_a_type;
  assign T_607 = T_606 ? 3'h3 : T_605;
  assign T_608 = 3'h1 == acq_io_deq_bits_a_type;
  assign T_609 = T_608 ? 3'h5 : T_607;
  assign T_610 = 3'h0 == acq_io_deq_bits_a_type;
  assign T_611 = T_610 ? 3'h4 : T_609;
  assign T_636_addr_beat = 3'h0;
  assign T_636_client_xact_id = acq_io_deq_bits_client_xact_id;
  assign T_636_manager_xact_id = 1'h0;
  assign T_636_is_builtin_type = 1'h1;
  assign T_636_g_type = {{1'd0}, T_611};
  assign T_636_data = rdata;
  assign T_658 = addr[15];
  assign T_660 = time$ + 64'h0;
  assign T_661 = T_660[63:0];
  assign T_667_0 = T_661;
  assign T_676_0 = 3'h0;
  assign T_676_1 = 3'h4;
  assign GEN_4 = T_658 ? T_667_0 : 64'h0;
  assign T_688 = addr >= 16'h4000;
  assign T_690 = T_658 == 1'h0;
  assign T_691 = T_690 & T_688;
  assign T_699_0 = 3'h0;
  assign T_699_1 = 3'h4;
  assign T_717_0 = 3'h0;
  assign T_717_1 = 3'h4;
  assign T_729 = acq_io_deq_bits_a_type == 3'h4;
  assign T_730 = acq_io_deq_bits_is_builtin_type & T_729;
  assign T_732 = T_574[2];
  assign T_734 = 2'h1 << T_732;
  assign T_735 = T_734[0];
  assign T_736 = T_734[1];
  assign T_740 = T_735 ? 4'hf : 4'h0;
  assign T_744 = T_736 ? 4'hf : 4'h0;
  assign T_745 = {T_744,T_740};
  assign T_747 = acq_io_deq_bits_a_type == 3'h3;
  assign T_748 = acq_io_deq_bits_is_builtin_type & T_747;
  assign T_750 = acq_io_deq_bits_a_type == 3'h2;
  assign T_751 = acq_io_deq_bits_is_builtin_type & T_750;
  assign T_752 = T_748 | T_751;
  assign T_753 = acq_io_deq_bits_union[8:1];
  assign T_755 = T_752 ? T_753 : 8'h0;
  assign T_756 = T_730 ? T_745 : T_755;
  assign T_757 = T_756[0];
  assign T_758 = T_756[1];
  assign T_759 = T_756[2];
  assign T_760 = T_756[3];
  assign T_761 = T_756[4];
  assign T_762 = T_756[5];
  assign T_763 = T_756[6];
  assign T_764 = T_756[7];
  assign T_768 = T_757 ? 8'hff : 8'h0;
  assign T_772 = T_758 ? 8'hff : 8'h0;
  assign T_776 = T_759 ? 8'hff : 8'h0;
  assign T_780 = T_760 ? 8'hff : 8'h0;
  assign T_784 = T_761 ? 8'hff : 8'h0;
  assign T_788 = T_762 ? 8'hff : 8'h0;
  assign T_792 = T_763 ? 8'hff : 8'h0;
  assign T_796 = T_764 ? 8'hff : 8'h0;
  assign T_797 = {T_772,T_768};
  assign T_798 = {T_780,T_776};
  assign T_799 = {T_798,T_797};
  assign T_800 = {T_788,T_784};
  assign T_801 = {T_796,T_792};
  assign T_802 = {T_801,T_800};
  assign T_803 = {T_802,T_799};
  assign T_804 = acq_io_deq_bits_data & T_803;
  assign T_881 = ~ T_803;
  assign T_882 = timecmp_0 & T_881;
  assign T_883 = T_804 | T_882;
  assign GEN_5 = T_751 ? T_883 : timecmp_0;
  assign GEN_10 = T_691 ? GEN_5 : timecmp_0;
  assign GEN_11 = T_691 ? timecmp_0 : GEN_4;
  assign T_895 = T_688 == 1'h0;
  assign T_896 = T_690 & T_895;
  assign T_904_0 = 3'h0;
  assign T_904_1 = 3'h4;
  assign T_922_0 = 3'h0;
  assign T_922_1 = 3'h4;
  assign GEN_19 = {{32'd0}, ipi_0};
  assign T_1087 = GEN_19 & T_881;
  assign T_1088 = T_804 | T_1087;
  assign GEN_12 = T_751 ? T_1088 : {{32'd0}, ipi_0};
  assign T_1099 = GEN_19 & 64'h100000001;
  assign GEN_17 = T_896 ? GEN_12 : {{32'd0}, ipi_0};
  assign GEN_18 = T_896 ? T_1099 : GEN_11;
  assign T_1100 = ipi_0[0];
  assign T_1101 = time$ >= timecmp_0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_2 = {2{$random}};
  timecmp_0 = GEN_2[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_3 = {2{$random}};
  time$ = GEN_3[63:0];
  `endif
  `ifdef RANDOMIZE
  GEN_6 = {1{$random}};
  ipi_0 = GEN_6[31:0];
  `endif
  `ifdef RANDOMIZE
  GEN_7 = {1{$random}};
  GEN_1 = GEN_7[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_691) begin
        if(T_751) begin
          timecmp_0 <= T_883;
        end
      end
    end
    if(reset) begin
      time$ <= 64'h0;
    end else begin
      if(io_rtcTick) begin
        time$ <= T_526;
      end
    end
    if(reset) begin
      ipi_0 <= T_533_0;
    end else begin
      ipi_0 <= GEN_17[31:0];
    end
  end
endmodule
module ROMSlave(
  input   clk,
  input   reset,
  output  io_acquire_ready,
  input   io_acquire_valid,
  input  [25:0] io_acquire_bits_addr_block,
  input  [1:0] io_acquire_bits_client_xact_id,
  input  [2:0] io_acquire_bits_addr_beat,
  input   io_acquire_bits_is_builtin_type,
  input  [2:0] io_acquire_bits_a_type,
  input  [11:0] io_acquire_bits_union,
  input  [63:0] io_acquire_bits_data,
  input   io_grant_ready,
  output  io_grant_valid,
  output [2:0] io_grant_bits_addr_beat,
  output [1:0] io_grant_bits_client_xact_id,
  output  io_grant_bits_manager_xact_id,
  output  io_grant_bits_is_builtin_type,
  output [3:0] io_grant_bits_g_type,
  output [63:0] io_grant_bits_data
);
  wire  acq_clk;
  wire  acq_reset;
  wire  acq_io_enq_ready;
  wire  acq_io_enq_valid;
  wire [25:0] acq_io_enq_bits_addr_block;
  wire [1:0] acq_io_enq_bits_client_xact_id;
  wire [2:0] acq_io_enq_bits_addr_beat;
  wire  acq_io_enq_bits_is_builtin_type;
  wire [2:0] acq_io_enq_bits_a_type;
  wire [11:0] acq_io_enq_bits_union;
  wire [63:0] acq_io_enq_bits_data;
  wire  acq_io_deq_ready;
  wire  acq_io_deq_valid;
  wire [25:0] acq_io_deq_bits_addr_block;
  wire [1:0] acq_io_deq_bits_client_xact_id;
  wire [2:0] acq_io_deq_bits_addr_beat;
  wire  acq_io_deq_bits_is_builtin_type;
  wire [2:0] acq_io_deq_bits_a_type;
  wire [11:0] acq_io_deq_bits_union;
  wire [63:0] acq_io_deq_bits_data;
  wire  acq_io_count;
  wire  T_446;
  wire  single_beat;
  wire  T_448;
  wire  multi_beat;
  wire  T_450;
  wire  T_451;
  wire  T_452;
  wire  T_453;
  wire  T_455;
  reg [2:0] addr_beat;
  reg [31:0] GEN_54;
  wire  T_457;
  wire [3:0] T_459;
  wire [2:0] T_460;
  wire [2:0] GEN_1;
  wire  T_461;
  wire [2:0] GEN_2;
  wire [63:0] rom_0;
  wire [63:0] rom_1;
  wire [63:0] rom_2;
  wire [63:0] rom_3;
  wire [63:0] rom_4;
  wire [63:0] rom_5;
  wire [63:0] rom_6;
  wire [63:0] rom_7;
  wire [63:0] rom_8;
  wire [63:0] rom_9;
  wire [63:0] rom_10;
  wire [63:0] rom_11;
  wire [63:0] rom_12;
  wire [63:0] rom_13;
  wire [63:0] rom_14;
  wire [63:0] rom_15;
  wire [63:0] rom_16;
  wire [63:0] rom_17;
  wire [63:0] rom_18;
  wire [63:0] rom_19;
  wire [63:0] rom_20;
  wire [63:0] rom_21;
  wire [63:0] rom_22;
  wire [63:0] rom_23;
  wire [63:0] rom_24;
  wire [63:0] rom_25;
  wire [63:0] rom_26;
  wire [63:0] rom_27;
  wire [63:0] rom_28;
  wire [63:0] rom_29;
  wire [63:0] rom_30;
  wire [63:0] rom_31;
  wire [63:0] rom_32;
  wire [63:0] rom_33;
  wire [63:0] rom_34;
  wire [63:0] rom_35;
  wire [63:0] rom_36;
  wire [63:0] rom_37;
  wire [63:0] rom_38;
  wire [63:0] rom_39;
  wire [63:0] rom_40;
  wire [63:0] rom_41;
  wire [63:0] rom_42;
  wire [63:0] rom_43;
  wire [63:0] rom_44;
  wire [63:0] rom_45;
  wire [63:0] rom_46;
  wire [63:0] rom_47;
  wire [63:0] rom_48;
  wire [63:0] rom_49;
  wire [63:0] rom_50;
  wire [63:0] rom_51;
  wire [28:0] raddr;
  wire [5:0] T_520;
  wire  T_522;
  wire  T_524;
  wire  last;
  wire  T_525;
  wire  T_542;
  wire [2:0] T_543;
  wire  T_544;
  wire [2:0] T_545;
  wire  T_546;
  wire [2:0] T_547;
  wire  T_548;
  wire [2:0] T_549;
  wire  T_550;
  wire [2:0] T_551;
  wire  T_552;
  wire [2:0] T_553;
  wire  T_554;
  wire [2:0] T_555;
  wire [2:0] T_579_addr_beat;
  wire [1:0] T_579_client_xact_id;
  wire  T_579_manager_xact_id;
  wire  T_579_is_builtin_type;
  wire [3:0] T_579_g_type;
  wire [63:0] T_579_data;
  wire [63:0] GEN_0;
  wire [63:0] GEN_3;
  wire [63:0] GEN_4;
  wire [63:0] GEN_5;
  wire [63:0] GEN_6;
  wire [63:0] GEN_7;
  wire [63:0] GEN_8;
  wire [63:0] GEN_9;
  wire [63:0] GEN_10;
  wire [63:0] GEN_11;
  wire [63:0] GEN_12;
  wire [63:0] GEN_13;
  wire [63:0] GEN_14;
  wire [63:0] GEN_15;
  wire [63:0] GEN_16;
  wire [63:0] GEN_17;
  wire [63:0] GEN_18;
  wire [63:0] GEN_19;
  wire [63:0] GEN_20;
  wire [63:0] GEN_21;
  wire [63:0] GEN_22;
  wire [63:0] GEN_23;
  wire [63:0] GEN_24;
  wire [63:0] GEN_25;
  wire [63:0] GEN_26;
  wire [63:0] GEN_27;
  wire [63:0] GEN_28;
  wire [63:0] GEN_29;
  wire [63:0] GEN_30;
  wire [63:0] GEN_31;
  wire [63:0] GEN_32;
  wire [63:0] GEN_33;
  wire [63:0] GEN_34;
  wire [63:0] GEN_35;
  wire [63:0] GEN_36;
  wire [63:0] GEN_37;
  wire [63:0] GEN_38;
  wire [63:0] GEN_39;
  wire [63:0] GEN_40;
  wire [63:0] GEN_41;
  wire [63:0] GEN_42;
  wire [63:0] GEN_43;
  wire [63:0] GEN_44;
  wire [63:0] GEN_45;
  wire [63:0] GEN_46;
  wire [63:0] GEN_47;
  wire [63:0] GEN_48;
  wire [63:0] GEN_49;
  wire [63:0] GEN_50;
  wire [63:0] GEN_51;
  wire [63:0] GEN_52;
  wire [63:0] GEN_53;
  Queue_8 acq (
    .clk(acq_clk),
    .reset(acq_reset),
    .io_enq_ready(acq_io_enq_ready),
    .io_enq_valid(acq_io_enq_valid),
    .io_enq_bits_addr_block(acq_io_enq_bits_addr_block),
    .io_enq_bits_client_xact_id(acq_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(acq_io_enq_bits_addr_beat),
    .io_enq_bits_is_builtin_type(acq_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(acq_io_enq_bits_a_type),
    .io_enq_bits_union(acq_io_enq_bits_union),
    .io_enq_bits_data(acq_io_enq_bits_data),
    .io_deq_ready(acq_io_deq_ready),
    .io_deq_valid(acq_io_deq_valid),
    .io_deq_bits_addr_block(acq_io_deq_bits_addr_block),
    .io_deq_bits_client_xact_id(acq_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(acq_io_deq_bits_addr_beat),
    .io_deq_bits_is_builtin_type(acq_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(acq_io_deq_bits_a_type),
    .io_deq_bits_union(acq_io_deq_bits_union),
    .io_deq_bits_data(acq_io_deq_bits_data),
    .io_count(acq_io_count)
  );
  assign io_acquire_ready = acq_io_enq_ready;
  assign io_grant_valid = acq_io_deq_valid;
  assign io_grant_bits_addr_beat = T_579_addr_beat;
  assign io_grant_bits_client_xact_id = T_579_client_xact_id;
  assign io_grant_bits_manager_xact_id = T_579_manager_xact_id;
  assign io_grant_bits_is_builtin_type = T_579_is_builtin_type;
  assign io_grant_bits_g_type = T_579_g_type;
  assign io_grant_bits_data = T_579_data;
  assign acq_clk = clk;
  assign acq_reset = reset;
  assign acq_io_enq_valid = io_acquire_valid;
  assign acq_io_enq_bits_addr_block = io_acquire_bits_addr_block;
  assign acq_io_enq_bits_client_xact_id = io_acquire_bits_client_xact_id;
  assign acq_io_enq_bits_addr_beat = io_acquire_bits_addr_beat;
  assign acq_io_enq_bits_is_builtin_type = io_acquire_bits_is_builtin_type;
  assign acq_io_enq_bits_a_type = io_acquire_bits_a_type;
  assign acq_io_enq_bits_union = io_acquire_bits_union;
  assign acq_io_enq_bits_data = io_acquire_bits_data;
  assign acq_io_deq_ready = T_525;
  assign T_446 = acq_io_deq_bits_a_type == 3'h0;
  assign single_beat = acq_io_deq_bits_is_builtin_type & T_446;
  assign T_448 = acq_io_deq_bits_a_type == 3'h1;
  assign multi_beat = acq_io_deq_bits_is_builtin_type & T_448;
  assign T_450 = acq_io_deq_valid == 1'h0;
  assign T_451 = T_450 | single_beat;
  assign T_452 = T_451 | multi_beat;
  assign T_453 = T_452 | reset;
  assign T_455 = T_453 == 1'h0;
  assign T_457 = io_grant_ready & io_grant_valid;
  assign T_459 = addr_beat + 3'h1;
  assign T_460 = T_459[2:0];
  assign GEN_1 = T_457 ? T_460 : addr_beat;
  assign T_461 = io_acquire_ready & io_acquire_valid;
  assign GEN_2 = T_461 ? io_acquire_bits_addr_beat : GEN_1;
  assign rom_0 = 64'h6f;
  assign rom_1 = 64'h6000002000000000;
  assign rom_2 = 64'h0;
  assign rom_3 = 64'h0;
  assign rom_4 = 64'h200a7b2063696c70;
  assign rom_5 = 64'h7469726f69727020;
  assign rom_6 = 64'h3030303478302079;
  assign rom_7 = 64'h20200a3b30303030;
  assign rom_8 = 64'h20676e69646e6570;
  assign rom_9 = 64'h3031303030347830;
  assign rom_10 = 64'h646e20200a3b3030;
  assign rom_11 = 64'ha3b313320737665;
  assign rom_12 = 64'h7b206374720a3b7d;
  assign rom_13 = 64'h207264646120200a;
  assign rom_14 = 64'h6662303034347830;
  assign rom_15 = 64'h720a3b7d0a3b3866;
  assign rom_16 = 64'h3020200a7b206d61;
  assign rom_17 = 64'h61202020200a7b20;
  assign rom_18 = 64'h3038783020726464;
  assign rom_19 = 64'ha3b303030303030;
  assign rom_20 = 64'h657a697320202020;
  assign rom_21 = 64'h3030303031783020;
  assign rom_22 = 64'h7d20200a3b303030;
  assign rom_23 = 64'h726f630a3b7d0a3b;
  assign rom_24 = 64'h203020200a7b2065;
  assign rom_25 = 64'h2030202020200a7b;
  assign rom_26 = 64'h2020202020200a7b;
  assign rom_27 = 64'h3233767220617369;
  assign rom_28 = 64'h202020200a3b6d69;
  assign rom_29 = 64'h6d63656d69742020;
  assign rom_30 = 64'h3030343478302070;
  assign rom_31 = 64'h20200a3b30303034;
  assign rom_32 = 64'h2069706920202020;
  assign rom_33 = 64'h3030303034347830;
  assign rom_34 = 64'h202020200a3b3030;
  assign rom_35 = 64'h7b2063696c702020;
  assign rom_36 = 64'h202020202020200a;
  assign rom_37 = 64'h2020200a7b206d20;
  assign rom_38 = 64'h6569202020202020;
  assign rom_39 = 64'h3230303034783020;
  assign rom_40 = 64'h2020200a3b303030;
  assign rom_41 = 64'h6874202020202020;
  assign rom_42 = 64'h3478302068736572;
  assign rom_43 = 64'h3b30303030303230;
  assign rom_44 = 64'h202020202020200a;
  assign rom_45 = 64'h206d69616c632020;
  assign rom_46 = 64'h3030303230347830;
  assign rom_47 = 64'h202020200a3b3430;
  assign rom_48 = 64'h200a3b7d20202020;
  assign rom_49 = 64'ha3b7d2020202020;
  assign rom_50 = 64'h200a3b7d20202020;
  assign rom_51 = 64'ha3b7d0a3b7d20;
  assign raddr = {acq_io_deq_bits_addr_block,addr_beat};
  assign T_520 = raddr[5:0];
  assign T_522 = multi_beat == 1'h0;
  assign T_524 = addr_beat == 3'h7;
  assign last = T_522 | T_524;
  assign T_525 = io_grant_ready & last;
  assign T_542 = 3'h6 == acq_io_deq_bits_a_type;
  assign T_543 = T_542 ? 3'h1 : 3'h3;
  assign T_544 = 3'h5 == acq_io_deq_bits_a_type;
  assign T_545 = T_544 ? 3'h1 : T_543;
  assign T_546 = 3'h4 == acq_io_deq_bits_a_type;
  assign T_547 = T_546 ? 3'h4 : T_545;
  assign T_548 = 3'h3 == acq_io_deq_bits_a_type;
  assign T_549 = T_548 ? 3'h3 : T_547;
  assign T_550 = 3'h2 == acq_io_deq_bits_a_type;
  assign T_551 = T_550 ? 3'h3 : T_549;
  assign T_552 = 3'h1 == acq_io_deq_bits_a_type;
  assign T_553 = T_552 ? 3'h5 : T_551;
  assign T_554 = 3'h0 == acq_io_deq_bits_a_type;
  assign T_555 = T_554 ? 3'h4 : T_553;
  assign T_579_addr_beat = addr_beat;
  assign T_579_client_xact_id = acq_io_deq_bits_client_xact_id;
  assign T_579_manager_xact_id = 1'h0;
  assign T_579_is_builtin_type = 1'h1;
  assign T_579_g_type = {{1'd0}, T_555};
  assign T_579_data = GEN_0;
  assign GEN_0 = GEN_53;
  assign GEN_3 = 6'h1 == T_520 ? rom_1 : rom_0;
  assign GEN_4 = 6'h2 == T_520 ? rom_2 : GEN_3;
  assign GEN_5 = 6'h3 == T_520 ? rom_3 : GEN_4;
  assign GEN_6 = 6'h4 == T_520 ? rom_4 : GEN_5;
  assign GEN_7 = 6'h5 == T_520 ? rom_5 : GEN_6;
  assign GEN_8 = 6'h6 == T_520 ? rom_6 : GEN_7;
  assign GEN_9 = 6'h7 == T_520 ? rom_7 : GEN_8;
  assign GEN_10 = 6'h8 == T_520 ? rom_8 : GEN_9;
  assign GEN_11 = 6'h9 == T_520 ? rom_9 : GEN_10;
  assign GEN_12 = 6'ha == T_520 ? rom_10 : GEN_11;
  assign GEN_13 = 6'hb == T_520 ? rom_11 : GEN_12;
  assign GEN_14 = 6'hc == T_520 ? rom_12 : GEN_13;
  assign GEN_15 = 6'hd == T_520 ? rom_13 : GEN_14;
  assign GEN_16 = 6'he == T_520 ? rom_14 : GEN_15;
  assign GEN_17 = 6'hf == T_520 ? rom_15 : GEN_16;
  assign GEN_18 = 6'h10 == T_520 ? rom_16 : GEN_17;
  assign GEN_19 = 6'h11 == T_520 ? rom_17 : GEN_18;
  assign GEN_20 = 6'h12 == T_520 ? rom_18 : GEN_19;
  assign GEN_21 = 6'h13 == T_520 ? rom_19 : GEN_20;
  assign GEN_22 = 6'h14 == T_520 ? rom_20 : GEN_21;
  assign GEN_23 = 6'h15 == T_520 ? rom_21 : GEN_22;
  assign GEN_24 = 6'h16 == T_520 ? rom_22 : GEN_23;
  assign GEN_25 = 6'h17 == T_520 ? rom_23 : GEN_24;
  assign GEN_26 = 6'h18 == T_520 ? rom_24 : GEN_25;
  assign GEN_27 = 6'h19 == T_520 ? rom_25 : GEN_26;
  assign GEN_28 = 6'h1a == T_520 ? rom_26 : GEN_27;
  assign GEN_29 = 6'h1b == T_520 ? rom_27 : GEN_28;
  assign GEN_30 = 6'h1c == T_520 ? rom_28 : GEN_29;
  assign GEN_31 = 6'h1d == T_520 ? rom_29 : GEN_30;
  assign GEN_32 = 6'h1e == T_520 ? rom_30 : GEN_31;
  assign GEN_33 = 6'h1f == T_520 ? rom_31 : GEN_32;
  assign GEN_34 = 6'h20 == T_520 ? rom_32 : GEN_33;
  assign GEN_35 = 6'h21 == T_520 ? rom_33 : GEN_34;
  assign GEN_36 = 6'h22 == T_520 ? rom_34 : GEN_35;
  assign GEN_37 = 6'h23 == T_520 ? rom_35 : GEN_36;
  assign GEN_38 = 6'h24 == T_520 ? rom_36 : GEN_37;
  assign GEN_39 = 6'h25 == T_520 ? rom_37 : GEN_38;
  assign GEN_40 = 6'h26 == T_520 ? rom_38 : GEN_39;
  assign GEN_41 = 6'h27 == T_520 ? rom_39 : GEN_40;
  assign GEN_42 = 6'h28 == T_520 ? rom_40 : GEN_41;
  assign GEN_43 = 6'h29 == T_520 ? rom_41 : GEN_42;
  assign GEN_44 = 6'h2a == T_520 ? rom_42 : GEN_43;
  assign GEN_45 = 6'h2b == T_520 ? rom_43 : GEN_44;
  assign GEN_46 = 6'h2c == T_520 ? rom_44 : GEN_45;
  assign GEN_47 = 6'h2d == T_520 ? rom_45 : GEN_46;
  assign GEN_48 = 6'h2e == T_520 ? rom_46 : GEN_47;
  assign GEN_49 = 6'h2f == T_520 ? rom_47 : GEN_48;
  assign GEN_50 = 6'h30 == T_520 ? rom_48 : GEN_49;
  assign GEN_51 = 6'h31 == T_520 ? rom_49 : GEN_50;
  assign GEN_52 = 6'h32 == T_520 ? rom_50 : GEN_51;
  assign GEN_53 = 6'h33 == T_520 ? rom_51 : GEN_52;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_54 = {1{$random}};
  addr_beat = GEN_54[2:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      if(T_461) begin
        addr_beat <= io_acquire_bits_addr_beat;
      end else begin
        if(T_457) begin
          addr_beat <= T_460;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_455) begin
          $fwrite(32'h80000002,"Assertion failed: unsupported ROMSlave operation\n    at Rom.scala:17 assert(!acq.valid || single_beat || multi_beat, ---unsupported ROMSlave operation---)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_455) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module ReorderQueue_3(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [2:0] io_enq_bits_data_addr_beat,
  input   io_enq_bits_data_subblock,
  input  [1:0] io_enq_bits_tag,
  input   io_deq_valid,
  input  [1:0] io_deq_tag,
  output [2:0] io_deq_data_addr_beat,
  output  io_deq_data_subblock,
  output  io_deq_matches
);
  reg [2:0] T_184_addr_beat [0:3];
  reg [31:0] GEN_14;
  wire [2:0] T_184_addr_beat_T_200_data;
  wire [1:0] T_184_addr_beat_T_200_addr;
  wire  T_184_addr_beat_T_200_en;
  wire [2:0] T_184_addr_beat_T_221_data;
  wire [1:0] T_184_addr_beat_T_221_addr;
  wire  T_184_addr_beat_T_221_mask;
  wire  T_184_addr_beat_T_221_en;
  reg  T_184_subblock [0:3];
  reg [31:0] GEN_15;
  wire  T_184_subblock_T_200_data;
  wire [1:0] T_184_subblock_T_200_addr;
  wire  T_184_subblock_T_200_en;
  wire  T_184_subblock_T_221_data;
  wire [1:0] T_184_subblock_T_221_addr;
  wire  T_184_subblock_T_221_mask;
  wire  T_184_subblock_T_221_en;
  wire  T_194_0;
  wire  T_194_1;
  wire  T_194_2;
  wire  T_194_3;
  reg  T_198_0;
  reg [31:0] GEN_16;
  reg  T_198_1;
  reg [31:0] GEN_17;
  reg  T_198_2;
  reg [31:0] GEN_18;
  reg  T_198_3;
  reg [31:0] GEN_19;
  wire  GEN_0;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_1;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  T_219;
  wire  T_220;
  wire  GEN_2;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_3;
  wire  GEN_26;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_29;
  wire  GEN_31;
  wire  GEN_32;
  wire  GEN_33;
  wire  GEN_34;
  assign io_enq_ready = GEN_0;
  assign io_deq_data_addr_beat = T_184_addr_beat_T_200_data;
  assign io_deq_data_subblock = T_184_subblock_T_200_data;
  assign io_deq_matches = T_219;
  assign T_184_addr_beat_T_200_addr = io_deq_tag;
  assign T_184_addr_beat_T_200_en = 1'h1;
  assign T_184_addr_beat_T_200_data = T_184_addr_beat[T_184_addr_beat_T_200_addr];
  assign T_184_addr_beat_T_221_data = io_enq_bits_data_addr_beat;
  assign T_184_addr_beat_T_221_addr = io_enq_bits_tag;
  assign T_184_addr_beat_T_221_mask = T_220;
  assign T_184_addr_beat_T_221_en = T_220;
  assign T_184_subblock_T_200_addr = io_deq_tag;
  assign T_184_subblock_T_200_en = 1'h1;
  assign T_184_subblock_T_200_data = T_184_subblock[T_184_subblock_T_200_addr];
  assign T_184_subblock_T_221_data = io_enq_bits_data_subblock;
  assign T_184_subblock_T_221_addr = io_enq_bits_tag;
  assign T_184_subblock_T_221_mask = T_220;
  assign T_184_subblock_T_221_en = T_220;
  assign T_194_0 = 1'h1;
  assign T_194_1 = 1'h1;
  assign T_194_2 = 1'h1;
  assign T_194_3 = 1'h1;
  assign GEN_0 = GEN_6;
  assign GEN_4 = 2'h1 == io_enq_bits_tag ? T_198_1 : T_198_0;
  assign GEN_5 = 2'h2 == io_enq_bits_tag ? T_198_2 : GEN_4;
  assign GEN_6 = 2'h3 == io_enq_bits_tag ? T_198_3 : GEN_5;
  assign GEN_1 = GEN_9;
  assign GEN_7 = 2'h1 == io_deq_tag ? T_198_1 : T_198_0;
  assign GEN_8 = 2'h2 == io_deq_tag ? T_198_2 : GEN_7;
  assign GEN_9 = 2'h3 == io_deq_tag ? T_198_3 : GEN_8;
  assign T_219 = GEN_1 == 1'h0;
  assign T_220 = io_enq_valid & io_enq_ready;
  assign GEN_2 = 1'h0;
  assign GEN_10 = 2'h0 == io_enq_bits_tag ? GEN_2 : T_198_0;
  assign GEN_11 = 2'h1 == io_enq_bits_tag ? GEN_2 : T_198_1;
  assign GEN_12 = 2'h2 == io_enq_bits_tag ? GEN_2 : T_198_2;
  assign GEN_13 = 2'h3 == io_enq_bits_tag ? GEN_2 : T_198_3;
  assign GEN_22 = T_220 ? GEN_10 : T_198_0;
  assign GEN_23 = T_220 ? GEN_11 : T_198_1;
  assign GEN_24 = T_220 ? GEN_12 : T_198_2;
  assign GEN_25 = T_220 ? GEN_13 : T_198_3;
  assign GEN_3 = 1'h1;
  assign GEN_26 = 2'h0 == io_deq_tag ? GEN_3 : GEN_22;
  assign GEN_27 = 2'h1 == io_deq_tag ? GEN_3 : GEN_23;
  assign GEN_28 = 2'h2 == io_deq_tag ? GEN_3 : GEN_24;
  assign GEN_29 = 2'h3 == io_deq_tag ? GEN_3 : GEN_25;
  assign GEN_31 = io_deq_valid ? GEN_26 : GEN_22;
  assign GEN_32 = io_deq_valid ? GEN_27 : GEN_23;
  assign GEN_33 = io_deq_valid ? GEN_28 : GEN_24;
  assign GEN_34 = io_deq_valid ? GEN_29 : GEN_25;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_14 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    T_184_addr_beat[initvar] = GEN_14[2:0];
  `endif
  GEN_15 = {1{$random}};
  `ifdef RANDOMIZE
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    T_184_subblock[initvar] = GEN_15[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_16 = {1{$random}};
  T_198_0 = GEN_16[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_17 = {1{$random}};
  T_198_1 = GEN_17[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_18 = {1{$random}};
  T_198_2 = GEN_18[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_19 = {1{$random}};
  T_198_3 = GEN_19[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(T_184_addr_beat_T_221_en & T_184_addr_beat_T_221_mask) begin
      T_184_addr_beat[T_184_addr_beat_T_221_addr] <= T_184_addr_beat_T_221_data;
    end
    if(T_184_subblock_T_221_en & T_184_subblock_T_221_mask) begin
      T_184_subblock[T_184_subblock_T_221_addr] <= T_184_subblock_T_221_data;
    end
    if(reset) begin
      T_198_0 <= T_194_0;
    end else begin
      if(io_deq_valid) begin
        if(2'h0 == io_deq_tag) begin
          T_198_0 <= GEN_3;
        end else begin
          if(T_220) begin
            if(2'h0 == io_enq_bits_tag) begin
              T_198_0 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_220) begin
          if(2'h0 == io_enq_bits_tag) begin
            T_198_0 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_198_1 <= T_194_1;
    end else begin
      if(io_deq_valid) begin
        if(2'h1 == io_deq_tag) begin
          T_198_1 <= GEN_3;
        end else begin
          if(T_220) begin
            if(2'h1 == io_enq_bits_tag) begin
              T_198_1 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_220) begin
          if(2'h1 == io_enq_bits_tag) begin
            T_198_1 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_198_2 <= T_194_2;
    end else begin
      if(io_deq_valid) begin
        if(2'h2 == io_deq_tag) begin
          T_198_2 <= GEN_3;
        end else begin
          if(T_220) begin
            if(2'h2 == io_enq_bits_tag) begin
              T_198_2 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_220) begin
          if(2'h2 == io_enq_bits_tag) begin
            T_198_2 <= GEN_2;
          end
        end
      end
    end
    if(reset) begin
      T_198_3 <= T_194_3;
    end else begin
      if(io_deq_valid) begin
        if(2'h3 == io_deq_tag) begin
          T_198_3 <= GEN_3;
        end else begin
          if(T_220) begin
            if(2'h3 == io_enq_bits_tag) begin
              T_198_3 <= GEN_2;
            end
          end
        end
      end else begin
        if(T_220) begin
          if(2'h3 == io_enq_bits_tag) begin
            T_198_3 <= GEN_2;
          end
        end
      end
    end
  end
endmodule
module LockingArbiter_1(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  input   io_in_0_bits_client_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [1:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_is_builtin_type,
  input  [3:0] io_in_1_bits_g_type,
  input  [63:0] io_in_1_bits_data,
  input   io_in_1_bits_client_id,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_out_bits_client_id,
  output  io_chosen
);
  wire  choice;
  wire  GEN_0;
  wire  GEN_8;
  wire [2:0] GEN_1;
  wire [2:0] GEN_9;
  wire [1:0] GEN_2;
  wire [1:0] GEN_10;
  wire  GEN_3;
  wire  GEN_11;
  wire  GEN_4;
  wire  GEN_12;
  wire [3:0] GEN_5;
  wire [3:0] GEN_13;
  wire [63:0] GEN_6;
  wire [63:0] GEN_14;
  wire  GEN_7;
  wire  GEN_15;
  reg [2:0] T_636;
  reg [31:0] GEN_21;
  reg  T_638;
  reg [31:0] GEN_22;
  wire  T_640;
  wire [2:0] T_648_0;
  wire [3:0] GEN_20;
  wire  T_650;
  wire  T_651;
  wire  T_652;
  wire  T_654;
  wire  T_655;
  wire [3:0] T_659;
  wire [2:0] T_660;
  wire  GEN_16;
  wire [2:0] GEN_17;
  wire  GEN_18;
  wire  T_663;
  wire  T_665;
  wire  T_666;
  wire  T_667;
  wire  T_670;
  wire  T_671;
  wire  GEN_19;
  assign io_in_0_ready = T_667;
  assign io_in_1_ready = T_671;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_beat = GEN_1;
  assign io_out_bits_client_xact_id = GEN_2;
  assign io_out_bits_manager_xact_id = GEN_3;
  assign io_out_bits_is_builtin_type = GEN_4;
  assign io_out_bits_g_type = GEN_5;
  assign io_out_bits_data = GEN_6;
  assign io_out_bits_client_id = GEN_7;
  assign io_chosen = GEN_18;
  assign choice = GEN_19;
  assign GEN_0 = GEN_8;
  assign GEN_8 = io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_1 = GEN_9;
  assign GEN_9 = io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_2 = GEN_10;
  assign GEN_10 = io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_3 = GEN_11;
  assign GEN_11 = io_chosen ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign GEN_4 = GEN_12;
  assign GEN_12 = io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_5 = GEN_13;
  assign GEN_13 = io_chosen ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign GEN_6 = GEN_14;
  assign GEN_14 = io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_7 = GEN_15;
  assign GEN_15 = io_chosen ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign T_640 = T_636 != 3'h0;
  assign T_648_0 = 3'h5;
  assign GEN_20 = {{1'd0}, T_648_0};
  assign T_650 = io_out_bits_g_type == GEN_20;
  assign T_651 = io_out_bits_g_type == 4'h0;
  assign T_652 = io_out_bits_is_builtin_type ? T_650 : T_651;
  assign T_654 = io_out_ready & io_out_valid;
  assign T_655 = T_654 & T_652;
  assign T_659 = T_636 + 3'h1;
  assign T_660 = T_659[2:0];
  assign GEN_16 = T_655 ? io_chosen : T_638;
  assign GEN_17 = T_655 ? T_660 : T_636;
  assign GEN_18 = T_640 ? T_638 : choice;
  assign T_663 = io_in_0_valid == 1'h0;
  assign T_665 = T_638 == 1'h0;
  assign T_666 = T_640 ? T_665 : 1'h1;
  assign T_667 = T_666 & io_out_ready;
  assign T_670 = T_640 ? T_638 : T_663;
  assign T_671 = T_670 & io_out_ready;
  assign GEN_19 = io_in_0_valid ? 1'h0 : 1'h1;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_21 = {1{$random}};
  T_636 = GEN_21[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_22 = {1{$random}};
  T_638 = GEN_22[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_636 <= 3'h0;
    end else begin
      if(T_655) begin
        T_636 <= T_660;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_655) begin
        T_638 <= io_chosen;
      end
    end
  end
endmodule
module NastiIOTileLinkIOConverter_1(
  input   clk,
  input   reset,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [11:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data,
  input   io_nasti_aw_ready,
  output  io_nasti_aw_valid,
  output [31:0] io_nasti_aw_bits_addr,
  output [7:0] io_nasti_aw_bits_len,
  output [2:0] io_nasti_aw_bits_size,
  output [1:0] io_nasti_aw_bits_burst,
  output  io_nasti_aw_bits_lock,
  output [3:0] io_nasti_aw_bits_cache,
  output [2:0] io_nasti_aw_bits_prot,
  output [3:0] io_nasti_aw_bits_qos,
  output [3:0] io_nasti_aw_bits_region,
  output [4:0] io_nasti_aw_bits_id,
  output  io_nasti_aw_bits_user,
  input   io_nasti_w_ready,
  output  io_nasti_w_valid,
  output [63:0] io_nasti_w_bits_data,
  output  io_nasti_w_bits_last,
  output [4:0] io_nasti_w_bits_id,
  output [7:0] io_nasti_w_bits_strb,
  output  io_nasti_w_bits_user,
  output  io_nasti_b_ready,
  input   io_nasti_b_valid,
  input  [1:0] io_nasti_b_bits_resp,
  input  [4:0] io_nasti_b_bits_id,
  input   io_nasti_b_bits_user,
  input   io_nasti_ar_ready,
  output  io_nasti_ar_valid,
  output [31:0] io_nasti_ar_bits_addr,
  output [7:0] io_nasti_ar_bits_len,
  output [2:0] io_nasti_ar_bits_size,
  output [1:0] io_nasti_ar_bits_burst,
  output  io_nasti_ar_bits_lock,
  output [3:0] io_nasti_ar_bits_cache,
  output [2:0] io_nasti_ar_bits_prot,
  output [3:0] io_nasti_ar_bits_qos,
  output [3:0] io_nasti_ar_bits_region,
  output [4:0] io_nasti_ar_bits_id,
  output  io_nasti_ar_bits_user,
  output  io_nasti_r_ready,
  input   io_nasti_r_valid,
  input  [1:0] io_nasti_r_bits_resp,
  input  [63:0] io_nasti_r_bits_data,
  input   io_nasti_r_bits_last,
  input  [4:0] io_nasti_r_bits_id,
  input   io_nasti_r_bits_user
);
  wire [2:0] T_593_0;
  wire [2:0] T_593_1;
  wire [2:0] T_593_2;
  wire  T_595;
  wire  T_596;
  wire  T_597;
  wire  T_598;
  wire  T_599;
  wire  has_data;
  wire [2:0] T_608_0;
  wire [2:0] T_608_1;
  wire [2:0] T_608_2;
  wire  T_610;
  wire  T_611;
  wire  T_612;
  wire  T_613;
  wire  T_614;
  wire  is_subblock;
  wire [2:0] T_623_0;
  wire  T_625;
  wire  is_multibeat;
  wire  T_626;
  wire  T_627;
  reg [2:0] tl_cnt_out;
  reg [31:0] GEN_11;
  wire  T_630;
  wire [3:0] T_632;
  wire [2:0] T_633;
  wire [2:0] GEN_0;
  wire  tl_wrap_out;
  wire  T_635;
  wire  get_valid;
  wire  put_valid;
  wire  roq_clk;
  wire  roq_reset;
  wire  roq_io_enq_ready;
  wire  roq_io_enq_valid;
  wire [2:0] roq_io_enq_bits_data_addr_beat;
  wire  roq_io_enq_bits_data_subblock;
  wire [1:0] roq_io_enq_bits_tag;
  wire  roq_io_deq_valid;
  wire [1:0] roq_io_deq_tag;
  wire [2:0] roq_io_deq_data_addr_beat;
  wire  roq_io_deq_data_subblock;
  wire  roq_io_deq_matches;
  wire  get_id_mapper_clk;
  wire  get_id_mapper_reset;
  wire  get_id_mapper_io_req_valid;
  wire  get_id_mapper_io_req_ready;
  wire [1:0] get_id_mapper_io_req_in_id;
  wire [4:0] get_id_mapper_io_req_out_id;
  wire  get_id_mapper_io_resp_valid;
  wire  get_id_mapper_io_resp_matches;
  wire [4:0] get_id_mapper_io_resp_out_id;
  wire [1:0] get_id_mapper_io_resp_in_id;
  wire  put_id_mapper_clk;
  wire  put_id_mapper_reset;
  wire  put_id_mapper_io_req_valid;
  wire  put_id_mapper_io_req_ready;
  wire [1:0] put_id_mapper_io_req_in_id;
  wire [4:0] put_id_mapper_io_req_out_id;
  wire  put_id_mapper_io_resp_valid;
  wire  put_id_mapper_io_resp_matches;
  wire [4:0] put_id_mapper_io_resp_out_id;
  wire [1:0] put_id_mapper_io_resp_in_id;
  wire  T_655;
  wire  put_id_mask;
  wire  T_657;
  wire  put_id_ready;
  reg  w_inflight;
  reg [31:0] GEN_12;
  reg [4:0] w_id;
  reg [31:0] GEN_13;
  wire  aw_ready;
  wire  T_660;
  wire  T_662;
  wire  T_663;
  reg [2:0] nasti_cnt_out;
  reg [31:0] GEN_14;
  wire  T_666;
  wire [3:0] T_668;
  wire [2:0] T_669;
  wire [2:0] GEN_1;
  wire  nasti_wrap_out;
  wire  T_670;
  wire  T_671;
  wire  T_673;
  wire  T_674;
  wire  T_675;
  wire  T_676;
  wire  T_678;
  wire  T_679;
  wire  T_680;
  wire  T_681;
  wire  T_682;
  wire  T_684;
  wire [2:0] T_692_0;
  wire [2:0] T_692_1;
  wire  T_694;
  wire  T_695;
  wire  T_696;
  wire  T_697;
  wire [2:0] T_698;
  wire [2:0] T_700;
  wire [28:0] T_701;
  wire [31:0] T_702;
  wire [2:0] T_703;
  wire  T_713;
  wire [2:0] T_714;
  wire  T_715;
  wire [2:0] T_716;
  wire  T_717;
  wire [2:0] T_718;
  wire  T_719;
  wire [2:0] T_720;
  wire  T_721;
  wire [2:0] T_722;
  wire  T_723;
  wire [2:0] T_724;
  wire  T_725;
  wire [2:0] T_726;
  wire  T_727;
  wire [2:0] T_728;
  wire [2:0] T_730;
  wire [2:0] T_733;
  wire [31:0] T_746_addr;
  wire [7:0] T_746_len;
  wire [2:0] T_746_size;
  wire [1:0] T_746_burst;
  wire  T_746_lock;
  wire [3:0] T_746_cache;
  wire [2:0] T_746_prot;
  wire [3:0] T_746_qos;
  wire [3:0] T_746_region;
  wire [4:0] T_746_id;
  wire  T_746_user;
  wire  T_765;
  wire  T_766;
  wire  T_768;
  wire [1:0] T_770;
  wire  T_771;
  wire  T_772;
  wire [3:0] T_776;
  wire [3:0] T_780;
  wire [7:0] T_781;
  wire  T_783;
  wire  T_784;
  wire  T_786;
  wire  T_787;
  wire  T_788;
  wire [7:0] T_789;
  wire [7:0] T_791;
  wire [7:0] T_792;
  wire [7:0] T_793;
  wire  T_794;
  wire  T_795;
  wire  T_796;
  wire  T_797;
  wire  T_798;
  wire  T_799;
  wire  T_800;
  wire  T_801;
  wire  T_802;
  wire  T_803;
  wire  T_804;
  wire  T_805;
  wire  T_806;
  wire  T_807;
  wire  T_814;
  wire [1:0] T_815;
  wire [1:0] T_817;
  wire  T_818;
  wire  T_819;
  wire  T_820;
  wire  T_821;
  wire  T_822;
  wire  T_823;
  wire  T_824;
  wire  T_825;
  wire [2:0] T_826;
  wire [1:0] T_828;
  wire  T_829;
  wire  T_830;
  wire  T_831;
  wire  T_832;
  wire  T_833;
  wire  T_834;
  wire  T_835;
  wire  T_836;
  wire  T_837;
  wire  T_838;
  wire  T_839;
  wire  T_840;
  wire  T_841;
  wire  T_842;
  wire  T_843;
  wire  T_844;
  wire  T_845;
  wire  T_846;
  wire [3:0] put_offset;
  wire [1:0] put_size;
  wire  T_849;
  wire  T_850;
  wire  T_851;
  wire  T_852;
  wire [2:0] T_860_0;
  wire [2:0] T_860_1;
  wire  T_862;
  wire  T_863;
  wire  T_864;
  wire  T_865;
  wire [2:0] T_868;
  wire [31:0] T_870;
  wire [3:0] T_872;
  wire [31:0] GEN_7;
  wire [31:0] T_873;
  wire [1:0] T_875;
  wire [2:0] T_878;
  wire [31:0] T_891_addr;
  wire [7:0] T_891_len;
  wire [2:0] T_891_size;
  wire [1:0] T_891_burst;
  wire  T_891_lock;
  wire [3:0] T_891_cache;
  wire [2:0] T_891_prot;
  wire [3:0] T_891_qos;
  wire [3:0] T_891_region;
  wire [4:0] T_891_id;
  wire  T_891_user;
  wire  T_910;
  wire  T_943;
  wire  T_944;
  wire [63:0] T_951_data;
  wire  T_951_last;
  wire [4:0] T_951_id;
  wire [7:0] T_951_strb;
  wire  T_951_user;
  wire  T_958;
  wire  T_959;
  wire  T_960;
  wire  T_961;
  wire  T_962;
  wire  T_966;
  wire  T_967;
  wire  GEN_2;
  wire [4:0] GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire  T_970;
  wire [2:0] T_978_0;
  wire [3:0] GEN_8;
  wire  T_980;
  wire  T_981;
  wire  T_982;
  wire  T_984;
  reg [2:0] tl_cnt_in;
  reg [31:0] GEN_15;
  wire [3:0] T_989;
  wire [2:0] T_990;
  wire [2:0] GEN_6;
  wire  gnt_arb_clk;
  wire  gnt_arb_reset;
  wire  gnt_arb_io_in_0_ready;
  wire  gnt_arb_io_in_0_valid;
  wire [2:0] gnt_arb_io_in_0_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_0_bits_client_xact_id;
  wire  gnt_arb_io_in_0_bits_manager_xact_id;
  wire  gnt_arb_io_in_0_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_0_bits_g_type;
  wire [63:0] gnt_arb_io_in_0_bits_data;
  wire  gnt_arb_io_in_0_bits_client_id;
  wire  gnt_arb_io_in_1_ready;
  wire  gnt_arb_io_in_1_valid;
  wire [2:0] gnt_arb_io_in_1_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_1_bits_client_xact_id;
  wire  gnt_arb_io_in_1_bits_manager_xact_id;
  wire  gnt_arb_io_in_1_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_1_bits_g_type;
  wire [63:0] gnt_arb_io_in_1_bits_data;
  wire  gnt_arb_io_in_1_bits_client_id;
  wire  gnt_arb_io_out_ready;
  wire  gnt_arb_io_out_valid;
  wire [2:0] gnt_arb_io_out_bits_addr_beat;
  wire [1:0] gnt_arb_io_out_bits_client_xact_id;
  wire  gnt_arb_io_out_bits_manager_xact_id;
  wire  gnt_arb_io_out_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_out_bits_g_type;
  wire [63:0] gnt_arb_io_out_bits_data;
  wire  gnt_arb_io_out_bits_client_id;
  wire  gnt_arb_io_chosen;
  wire [2:0] T_1017;
  wire [2:0] T_1019;
  wire [2:0] T_1042_addr_beat;
  wire [1:0] T_1042_client_xact_id;
  wire  T_1042_manager_xact_id;
  wire  T_1042_is_builtin_type;
  wire [3:0] T_1042_g_type;
  wire [63:0] T_1042_data;
  wire  T_1065;
  wire  T_1066;
  wire  T_1067;
  wire  T_1069;
  wire  T_1071;
  wire  T_1072;
  wire  T_1073;
  wire  T_1075;
  wire [2:0] T_1103_addr_beat;
  wire [1:0] T_1103_client_xact_id;
  wire  T_1103_manager_xact_id;
  wire  T_1103_is_builtin_type;
  wire [3:0] T_1103_g_type;
  wire [63:0] T_1103_data;
  wire  T_1126;
  wire  T_1127;
  wire  T_1128;
  wire  T_1130;
  wire  T_1132;
  wire  T_1134;
  wire  T_1135;
  wire  T_1136;
  wire  T_1138;
  wire  T_1140;
  wire  T_1142;
  wire  T_1143;
  wire  T_1144;
  wire  T_1146;
  reg  GEN_9;
  reg [31:0] GEN_16;
  reg  GEN_10;
  reg [31:0] GEN_17;
  ReorderQueue_3 roq (
    .clk(roq_clk),
    .reset(roq_reset),
    .io_enq_ready(roq_io_enq_ready),
    .io_enq_valid(roq_io_enq_valid),
    .io_enq_bits_data_addr_beat(roq_io_enq_bits_data_addr_beat),
    .io_enq_bits_data_subblock(roq_io_enq_bits_data_subblock),
    .io_enq_bits_tag(roq_io_enq_bits_tag),
    .io_deq_valid(roq_io_deq_valid),
    .io_deq_tag(roq_io_deq_tag),
    .io_deq_data_addr_beat(roq_io_deq_data_addr_beat),
    .io_deq_data_subblock(roq_io_deq_data_subblock),
    .io_deq_matches(roq_io_deq_matches)
  );
  IdMapper get_id_mapper (
    .clk(get_id_mapper_clk),
    .reset(get_id_mapper_reset),
    .io_req_valid(get_id_mapper_io_req_valid),
    .io_req_ready(get_id_mapper_io_req_ready),
    .io_req_in_id(get_id_mapper_io_req_in_id),
    .io_req_out_id(get_id_mapper_io_req_out_id),
    .io_resp_valid(get_id_mapper_io_resp_valid),
    .io_resp_matches(get_id_mapper_io_resp_matches),
    .io_resp_out_id(get_id_mapper_io_resp_out_id),
    .io_resp_in_id(get_id_mapper_io_resp_in_id)
  );
  IdMapper put_id_mapper (
    .clk(put_id_mapper_clk),
    .reset(put_id_mapper_reset),
    .io_req_valid(put_id_mapper_io_req_valid),
    .io_req_ready(put_id_mapper_io_req_ready),
    .io_req_in_id(put_id_mapper_io_req_in_id),
    .io_req_out_id(put_id_mapper_io_req_out_id),
    .io_resp_valid(put_id_mapper_io_resp_valid),
    .io_resp_matches(put_id_mapper_io_resp_matches),
    .io_resp_out_id(put_id_mapper_io_resp_out_id),
    .io_resp_in_id(put_id_mapper_io_resp_in_id)
  );
  LockingArbiter_1 gnt_arb (
    .clk(gnt_arb_clk),
    .reset(gnt_arb_reset),
    .io_in_0_ready(gnt_arb_io_in_0_ready),
    .io_in_0_valid(gnt_arb_io_in_0_valid),
    .io_in_0_bits_addr_beat(gnt_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(gnt_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(gnt_arb_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(gnt_arb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(gnt_arb_io_in_0_bits_g_type),
    .io_in_0_bits_data(gnt_arb_io_in_0_bits_data),
    .io_in_0_bits_client_id(gnt_arb_io_in_0_bits_client_id),
    .io_in_1_ready(gnt_arb_io_in_1_ready),
    .io_in_1_valid(gnt_arb_io_in_1_valid),
    .io_in_1_bits_addr_beat(gnt_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_client_xact_id(gnt_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_manager_xact_id(gnt_arb_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_is_builtin_type(gnt_arb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_g_type(gnt_arb_io_in_1_bits_g_type),
    .io_in_1_bits_data(gnt_arb_io_in_1_bits_data),
    .io_in_1_bits_client_id(gnt_arb_io_in_1_bits_client_id),
    .io_out_ready(gnt_arb_io_out_ready),
    .io_out_valid(gnt_arb_io_out_valid),
    .io_out_bits_addr_beat(gnt_arb_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(gnt_arb_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(gnt_arb_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(gnt_arb_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(gnt_arb_io_out_bits_g_type),
    .io_out_bits_data(gnt_arb_io_out_bits_data),
    .io_out_bits_client_id(gnt_arb_io_out_bits_client_id),
    .io_chosen(gnt_arb_io_chosen)
  );
  assign io_tl_acquire_ready = T_962;
  assign io_tl_grant_valid = gnt_arb_io_out_valid;
  assign io_tl_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_tl_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_tl_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_tl_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_nasti_aw_valid = T_852;
  assign io_nasti_aw_bits_addr = T_891_addr;
  assign io_nasti_aw_bits_len = T_891_len;
  assign io_nasti_aw_bits_size = T_891_size;
  assign io_nasti_aw_bits_burst = T_891_burst;
  assign io_nasti_aw_bits_lock = T_891_lock;
  assign io_nasti_aw_bits_cache = T_891_cache;
  assign io_nasti_aw_bits_prot = T_891_prot;
  assign io_nasti_aw_bits_qos = T_891_qos;
  assign io_nasti_aw_bits_region = T_891_region;
  assign io_nasti_aw_bits_id = T_891_id;
  assign io_nasti_aw_bits_user = T_891_user;
  assign io_nasti_w_valid = T_910;
  assign io_nasti_w_bits_data = T_951_data;
  assign io_nasti_w_bits_last = T_951_last;
  assign io_nasti_w_bits_id = T_951_id;
  assign io_nasti_w_bits_strb = T_951_strb;
  assign io_nasti_w_bits_user = T_951_user;
  assign io_nasti_b_ready = gnt_arb_io_in_1_ready;
  assign io_nasti_ar_valid = T_684;
  assign io_nasti_ar_bits_addr = T_746_addr;
  assign io_nasti_ar_bits_len = T_746_len;
  assign io_nasti_ar_bits_size = T_746_size;
  assign io_nasti_ar_bits_burst = T_746_burst;
  assign io_nasti_ar_bits_lock = T_746_lock;
  assign io_nasti_ar_bits_cache = T_746_cache;
  assign io_nasti_ar_bits_prot = T_746_prot;
  assign io_nasti_ar_bits_qos = T_746_qos;
  assign io_nasti_ar_bits_region = T_746_region;
  assign io_nasti_ar_bits_id = T_746_id;
  assign io_nasti_ar_bits_user = T_746_user;
  assign io_nasti_r_ready = gnt_arb_io_in_0_ready;
  assign T_593_0 = 3'h2;
  assign T_593_1 = 3'h3;
  assign T_593_2 = 3'h4;
  assign T_595 = io_tl_acquire_bits_a_type == T_593_0;
  assign T_596 = io_tl_acquire_bits_a_type == T_593_1;
  assign T_597 = io_tl_acquire_bits_a_type == T_593_2;
  assign T_598 = T_595 | T_596;
  assign T_599 = T_598 | T_597;
  assign has_data = io_tl_acquire_bits_is_builtin_type & T_599;
  assign T_608_0 = 3'h2;
  assign T_608_1 = 3'h0;
  assign T_608_2 = 3'h4;
  assign T_610 = io_tl_acquire_bits_a_type == T_608_0;
  assign T_611 = io_tl_acquire_bits_a_type == T_608_1;
  assign T_612 = io_tl_acquire_bits_a_type == T_608_2;
  assign T_613 = T_610 | T_611;
  assign T_614 = T_613 | T_612;
  assign is_subblock = io_tl_acquire_bits_is_builtin_type & T_614;
  assign T_623_0 = 3'h3;
  assign T_625 = io_tl_acquire_bits_a_type == T_623_0;
  assign is_multibeat = io_tl_acquire_bits_is_builtin_type & T_625;
  assign T_626 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign T_627 = T_626 & is_multibeat;
  assign T_630 = tl_cnt_out == 3'h7;
  assign T_632 = tl_cnt_out + 3'h1;
  assign T_633 = T_632[2:0];
  assign GEN_0 = T_627 ? T_633 : tl_cnt_out;
  assign tl_wrap_out = T_627 & T_630;
  assign T_635 = has_data == 1'h0;
  assign get_valid = io_tl_acquire_valid & T_635;
  assign put_valid = io_tl_acquire_valid & has_data;
  assign roq_clk = clk;
  assign roq_reset = reset;
  assign roq_io_enq_valid = T_671;
  assign roq_io_enq_bits_data_addr_beat = io_tl_acquire_bits_addr_beat;
  assign roq_io_enq_bits_data_subblock = is_subblock;
  assign roq_io_enq_bits_tag = io_nasti_ar_bits_id[1:0];
  assign roq_io_deq_valid = T_674;
  assign roq_io_deq_tag = io_nasti_r_bits_id[1:0];
  assign get_id_mapper_clk = clk;
  assign get_id_mapper_reset = reset;
  assign get_id_mapper_io_req_valid = T_676;
  assign get_id_mapper_io_req_in_id = io_tl_acquire_bits_client_xact_id;
  assign get_id_mapper_io_resp_valid = T_678;
  assign get_id_mapper_io_resp_out_id = io_nasti_r_bits_id;
  assign put_id_mapper_clk = clk;
  assign put_id_mapper_reset = reset;
  assign put_id_mapper_io_req_valid = T_681;
  assign put_id_mapper_io_req_in_id = io_tl_acquire_bits_client_xact_id;
  assign put_id_mapper_io_resp_valid = T_682;
  assign put_id_mapper_io_resp_out_id = io_nasti_b_bits_id;
  assign T_655 = io_tl_acquire_bits_addr_beat == 3'h0;
  assign put_id_mask = is_subblock | T_655;
  assign T_657 = put_id_mask == 1'h0;
  assign put_id_ready = put_id_mapper_io_req_ready | T_657;
  assign aw_ready = w_inflight | io_nasti_aw_ready;
  assign T_660 = io_nasti_r_ready & io_nasti_r_valid;
  assign T_662 = roq_io_deq_data_subblock == 1'h0;
  assign T_663 = T_660 & T_662;
  assign T_666 = nasti_cnt_out == 3'h7;
  assign T_668 = nasti_cnt_out + 3'h1;
  assign T_669 = T_668[2:0];
  assign GEN_1 = T_663 ? T_669 : nasti_cnt_out;
  assign nasti_wrap_out = T_663 & T_666;
  assign T_670 = get_valid & io_nasti_ar_ready;
  assign T_671 = T_670 & get_id_mapper_io_req_ready;
  assign T_673 = nasti_wrap_out | roq_io_deq_data_subblock;
  assign T_674 = T_660 & T_673;
  assign T_675 = get_valid & roq_io_enq_ready;
  assign T_676 = T_675 & io_nasti_ar_ready;
  assign T_678 = T_660 & io_nasti_r_bits_last;
  assign T_679 = put_valid & aw_ready;
  assign T_680 = T_679 & io_nasti_w_ready;
  assign T_681 = T_680 & put_id_mask;
  assign T_682 = io_nasti_b_ready & io_nasti_b_valid;
  assign T_684 = T_675 & get_id_mapper_io_req_ready;
  assign T_692_0 = 3'h0;
  assign T_692_1 = 3'h4;
  assign T_694 = io_tl_acquire_bits_a_type == T_692_0;
  assign T_695 = io_tl_acquire_bits_a_type == T_692_1;
  assign T_696 = T_694 | T_695;
  assign T_697 = io_tl_acquire_bits_is_builtin_type & T_696;
  assign T_698 = io_tl_acquire_bits_union[11:9];
  assign T_700 = T_697 ? T_698 : 3'h0;
  assign T_701 = {io_tl_acquire_bits_addr_block,io_tl_acquire_bits_addr_beat};
  assign T_702 = {T_701,T_700};
  assign T_703 = io_tl_acquire_bits_union[8:6];
  assign T_713 = 3'h7 == T_703;
  assign T_714 = T_713 ? 3'h3 : 3'h7;
  assign T_715 = 3'h3 == T_703;
  assign T_716 = T_715 ? 3'h3 : T_714;
  assign T_717 = 3'h6 == T_703;
  assign T_718 = T_717 ? 3'h2 : T_716;
  assign T_719 = 3'h2 == T_703;
  assign T_720 = T_719 ? 3'h2 : T_718;
  assign T_721 = 3'h5 == T_703;
  assign T_722 = T_721 ? 3'h1 : T_720;
  assign T_723 = 3'h1 == T_703;
  assign T_724 = T_723 ? 3'h1 : T_722;
  assign T_725 = 3'h4 == T_703;
  assign T_726 = T_725 ? 3'h0 : T_724;
  assign T_727 = 3'h0 == T_703;
  assign T_728 = T_727 ? 3'h0 : T_726;
  assign T_730 = is_subblock ? T_728 : 3'h3;
  assign T_733 = is_subblock ? 3'h0 : 3'h7;
  assign T_746_addr = T_702;
  assign T_746_len = {{5'd0}, T_733};
  assign T_746_size = T_730;
  assign T_746_burst = 2'h1;
  assign T_746_lock = 1'h0;
  assign T_746_cache = 4'h0;
  assign T_746_prot = 3'h0;
  assign T_746_qos = 4'h0;
  assign T_746_region = 4'h0;
  assign T_746_id = get_id_mapper_io_req_out_id;
  assign T_746_user = 1'h0;
  assign T_765 = io_tl_acquire_bits_a_type == 3'h4;
  assign T_766 = io_tl_acquire_bits_is_builtin_type & T_765;
  assign T_768 = T_698[2];
  assign T_770 = 2'h1 << T_768;
  assign T_771 = T_770[0];
  assign T_772 = T_770[1];
  assign T_776 = T_771 ? 4'hf : 4'h0;
  assign T_780 = T_772 ? 4'hf : 4'h0;
  assign T_781 = {T_780,T_776};
  assign T_783 = io_tl_acquire_bits_a_type == 3'h3;
  assign T_784 = io_tl_acquire_bits_is_builtin_type & T_783;
  assign T_786 = io_tl_acquire_bits_a_type == 3'h2;
  assign T_787 = io_tl_acquire_bits_is_builtin_type & T_786;
  assign T_788 = T_784 | T_787;
  assign T_789 = io_tl_acquire_bits_union[8:1];
  assign T_791 = T_788 ? T_789 : 8'h0;
  assign T_792 = T_766 ? T_781 : T_791;
  assign T_793 = ~ T_792;
  assign T_794 = T_793[0];
  assign T_795 = T_793[1];
  assign T_796 = T_793[2];
  assign T_797 = T_793[3];
  assign T_798 = T_793[4];
  assign T_799 = T_793[5];
  assign T_800 = T_793[6];
  assign T_801 = T_793[7];
  assign T_802 = T_794 & T_795;
  assign T_803 = T_796 & T_797;
  assign T_804 = T_798 & T_799;
  assign T_805 = T_800 & T_801;
  assign T_806 = T_802 & T_803;
  assign T_807 = T_804 & T_805;
  assign T_814 = T_807 | T_806;
  assign T_815 = {1'h0,T_806};
  assign T_817 = T_814 ? 2'h2 : 2'h3;
  assign T_818 = T_807 & T_803;
  assign T_819 = T_807 & T_802;
  assign T_820 = T_806 & T_805;
  assign T_821 = T_806 & T_804;
  assign T_822 = T_819 | T_821;
  assign T_823 = T_818 | T_819;
  assign T_824 = T_823 | T_820;
  assign T_825 = T_824 | T_821;
  assign T_826 = {T_815,T_822};
  assign T_828 = T_825 ? 2'h1 : T_817;
  assign T_829 = T_818 & T_795;
  assign T_830 = T_818 & T_794;
  assign T_831 = T_819 & T_797;
  assign T_832 = T_819 & T_796;
  assign T_833 = T_820 & T_799;
  assign T_834 = T_820 & T_798;
  assign T_835 = T_821 & T_801;
  assign T_836 = T_821 & T_800;
  assign T_837 = T_830 | T_832;
  assign T_838 = T_837 | T_834;
  assign T_839 = T_838 | T_836;
  assign T_840 = T_829 | T_830;
  assign T_841 = T_840 | T_831;
  assign T_842 = T_841 | T_832;
  assign T_843 = T_842 | T_833;
  assign T_844 = T_843 | T_834;
  assign T_845 = T_844 | T_835;
  assign T_846 = T_845 | T_836;
  assign put_offset = {T_826,T_839};
  assign put_size = T_846 ? 2'h0 : T_828;
  assign T_849 = w_inflight == 1'h0;
  assign T_850 = put_valid & io_nasti_w_ready;
  assign T_851 = T_850 & put_id_ready;
  assign T_852 = T_851 & T_849;
  assign T_860_0 = 3'h0;
  assign T_860_1 = 3'h4;
  assign T_862 = io_tl_acquire_bits_a_type == T_860_0;
  assign T_863 = io_tl_acquire_bits_a_type == T_860_1;
  assign T_864 = T_862 | T_863;
  assign T_865 = io_tl_acquire_bits_is_builtin_type & T_864;
  assign T_868 = T_865 ? T_698 : 3'h0;
  assign T_870 = {T_701,T_868};
  assign T_872 = is_multibeat ? 4'h0 : put_offset;
  assign GEN_7 = {{28'd0}, T_872};
  assign T_873 = T_870 | GEN_7;
  assign T_875 = is_multibeat ? 2'h3 : put_size;
  assign T_878 = is_multibeat ? 3'h7 : 3'h0;
  assign T_891_addr = T_873;
  assign T_891_len = {{5'd0}, T_878};
  assign T_891_size = {{1'd0}, T_875};
  assign T_891_burst = 2'h1;
  assign T_891_lock = 1'h0;
  assign T_891_cache = 4'h0;
  assign T_891_prot = 3'h0;
  assign T_891_qos = 4'h0;
  assign T_891_region = 4'h0;
  assign T_891_id = put_id_mapper_io_req_out_id;
  assign T_891_user = 1'h0;
  assign T_910 = T_679 & put_id_ready;
  assign T_943 = is_multibeat == 1'h0;
  assign T_944 = w_inflight ? T_630 : T_943;
  assign T_951_data = io_tl_acquire_bits_data;
  assign T_951_last = T_944;
  assign T_951_id = w_id;
  assign T_951_strb = T_792;
  assign T_951_user = 1'h0;
  assign T_958 = aw_ready & io_nasti_w_ready;
  assign T_959 = T_958 & put_id_ready;
  assign T_960 = roq_io_enq_ready & io_nasti_ar_ready;
  assign T_961 = T_960 & get_id_mapper_io_req_ready;
  assign T_962 = has_data ? T_959 : T_961;
  assign T_966 = T_849 & T_626;
  assign T_967 = T_966 & is_multibeat;
  assign GEN_2 = T_967 ? 1'h1 : w_inflight;
  assign GEN_3 = T_967 ? put_id_mapper_io_req_out_id : w_id;
  assign GEN_4 = tl_wrap_out ? 1'h0 : GEN_2;
  assign GEN_5 = w_inflight ? GEN_4 : GEN_2;
  assign T_970 = io_tl_grant_ready & io_tl_grant_valid;
  assign T_978_0 = 3'h5;
  assign GEN_8 = {{1'd0}, T_978_0};
  assign T_980 = io_tl_grant_bits_g_type == GEN_8;
  assign T_981 = io_tl_grant_bits_g_type == 4'h0;
  assign T_982 = io_tl_grant_bits_is_builtin_type ? T_980 : T_981;
  assign T_984 = T_970 & T_982;
  assign T_989 = tl_cnt_in + 3'h1;
  assign T_990 = T_989[2:0];
  assign GEN_6 = T_984 ? T_990 : tl_cnt_in;
  assign gnt_arb_clk = clk;
  assign gnt_arb_reset = reset;
  assign gnt_arb_io_in_0_valid = io_nasti_r_valid;
  assign gnt_arb_io_in_0_bits_addr_beat = T_1042_addr_beat;
  assign gnt_arb_io_in_0_bits_client_xact_id = T_1042_client_xact_id;
  assign gnt_arb_io_in_0_bits_manager_xact_id = T_1042_manager_xact_id;
  assign gnt_arb_io_in_0_bits_is_builtin_type = T_1042_is_builtin_type;
  assign gnt_arb_io_in_0_bits_g_type = T_1042_g_type;
  assign gnt_arb_io_in_0_bits_data = T_1042_data;
  assign gnt_arb_io_in_0_bits_client_id = GEN_9;
  assign gnt_arb_io_in_1_valid = io_nasti_b_valid;
  assign gnt_arb_io_in_1_bits_addr_beat = T_1103_addr_beat;
  assign gnt_arb_io_in_1_bits_client_xact_id = T_1103_client_xact_id;
  assign gnt_arb_io_in_1_bits_manager_xact_id = T_1103_manager_xact_id;
  assign gnt_arb_io_in_1_bits_is_builtin_type = T_1103_is_builtin_type;
  assign gnt_arb_io_in_1_bits_g_type = T_1103_g_type;
  assign gnt_arb_io_in_1_bits_data = T_1103_data;
  assign gnt_arb_io_in_1_bits_client_id = GEN_10;
  assign gnt_arb_io_out_ready = io_tl_grant_ready;
  assign T_1017 = roq_io_deq_data_subblock ? 3'h4 : 3'h5;
  assign T_1019 = roq_io_deq_data_subblock ? roq_io_deq_data_addr_beat : tl_cnt_in;
  assign T_1042_addr_beat = T_1019;
  assign T_1042_client_xact_id = get_id_mapper_io_resp_in_id;
  assign T_1042_manager_xact_id = 1'h0;
  assign T_1042_is_builtin_type = 1'h1;
  assign T_1042_g_type = {{1'd0}, T_1017};
  assign T_1042_data = io_nasti_r_bits_data;
  assign T_1065 = roq_io_deq_valid == 1'h0;
  assign T_1066 = T_1065 | roq_io_deq_matches;
  assign T_1067 = T_1066 | reset;
  assign T_1069 = T_1067 == 1'h0;
  assign T_1071 = gnt_arb_io_in_0_valid == 1'h0;
  assign T_1072 = T_1071 | get_id_mapper_io_resp_matches;
  assign T_1073 = T_1072 | reset;
  assign T_1075 = T_1073 == 1'h0;
  assign T_1103_addr_beat = 3'h0;
  assign T_1103_client_xact_id = put_id_mapper_io_resp_in_id;
  assign T_1103_manager_xact_id = 1'h0;
  assign T_1103_is_builtin_type = 1'h1;
  assign T_1103_g_type = 4'h3;
  assign T_1103_data = 64'h0;
  assign T_1126 = gnt_arb_io_in_1_valid == 1'h0;
  assign T_1127 = T_1126 | put_id_mapper_io_resp_matches;
  assign T_1128 = T_1127 | reset;
  assign T_1130 = T_1128 == 1'h0;
  assign T_1132 = io_nasti_r_valid == 1'h0;
  assign T_1134 = io_nasti_r_bits_resp == 2'h0;
  assign T_1135 = T_1132 | T_1134;
  assign T_1136 = T_1135 | reset;
  assign T_1138 = T_1136 == 1'h0;
  assign T_1140 = io_nasti_b_valid == 1'h0;
  assign T_1142 = io_nasti_b_bits_resp == 2'h0;
  assign T_1143 = T_1140 | T_1142;
  assign T_1144 = T_1143 | reset;
  assign T_1146 = T_1144 == 1'h0;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_11 = {1{$random}};
  tl_cnt_out = GEN_11[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_12 = {1{$random}};
  w_inflight = GEN_12[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_13 = {1{$random}};
  w_id = GEN_13[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_14 = {1{$random}};
  nasti_cnt_out = GEN_14[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_15 = {1{$random}};
  tl_cnt_in = GEN_15[2:0];
  `endif
  `ifdef RANDOMIZE
  GEN_16 = {1{$random}};
  GEN_9 = GEN_16[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_17 = {1{$random}};
  GEN_10 = GEN_17[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      tl_cnt_out <= 3'h0;
    end else begin
      if(T_627) begin
        tl_cnt_out <= T_633;
      end
    end
    if(reset) begin
      w_inflight <= 1'h0;
    end else begin
      if(w_inflight) begin
        if(tl_wrap_out) begin
          w_inflight <= 1'h0;
        end else begin
          if(T_967) begin
            w_inflight <= 1'h1;
          end
        end
      end else begin
        if(T_967) begin
          w_inflight <= 1'h1;
        end
      end
    end
    if(reset) begin
      w_id <= 5'h0;
    end else begin
      if(T_967) begin
        w_id <= put_id_mapper_io_req_out_id;
      end
    end
    if(reset) begin
      nasti_cnt_out <= 3'h0;
    end else begin
      if(T_663) begin
        nasti_cnt_out <= T_669;
      end
    end
    if(reset) begin
      tl_cnt_in <= 3'h0;
    end else begin
      if(T_984) begin
        tl_cnt_in <= T_990;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1069) begin
          $fwrite(32'h80000002,"Assertion failed: TL -> NASTI converter ReorderQueue: NASTI tag error\n    at Nasti.scala:229 assert(!roq.io.deq.valid || roq.io.deq.matches,\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1069) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1075) begin
          $fwrite(32'h80000002,"Assertion failed: TL -> NASTI ID Mapper: NASTI tag error\n    at Nasti.scala:231 assert(!gnt_arb.io.in(0).valid || get_id_mapper.io.resp.matches,\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1075) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1130) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI tag error\n    at Nasti.scala:243 assert(!gnt_arb.io.in(1).valid || put_id_mapper.io.resp.matches, ---NASTI tag error---)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1130) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1138) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI read error\n    at Nasti.scala:245 assert(!io.nasti.r.valid || io.nasti.r.bits.resp === UInt(0), ---NASTI read error---)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1138) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1146) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI write error\n    at Nasti.scala:246 assert(!io.nasti.b.valid || io.nasti.b.bits.resp === UInt(0), ---NASTI write error---)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1146) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
module Uncore(
  input   clk,
  input   reset,
  input   io_mem_axi_0_aw_ready,
  output  io_mem_axi_0_aw_valid,
  output [31:0] io_mem_axi_0_aw_bits_addr,
  output [7:0] io_mem_axi_0_aw_bits_len,
  output [2:0] io_mem_axi_0_aw_bits_size,
  output [1:0] io_mem_axi_0_aw_bits_burst,
  output  io_mem_axi_0_aw_bits_lock,
  output [3:0] io_mem_axi_0_aw_bits_cache,
  output [2:0] io_mem_axi_0_aw_bits_prot,
  output [3:0] io_mem_axi_0_aw_bits_qos,
  output [3:0] io_mem_axi_0_aw_bits_region,
  output [4:0] io_mem_axi_0_aw_bits_id,
  output  io_mem_axi_0_aw_bits_user,
  input   io_mem_axi_0_w_ready,
  output  io_mem_axi_0_w_valid,
  output [63:0] io_mem_axi_0_w_bits_data,
  output  io_mem_axi_0_w_bits_last,
  output [4:0] io_mem_axi_0_w_bits_id,
  output [7:0] io_mem_axi_0_w_bits_strb,
  output  io_mem_axi_0_w_bits_user,
  output  io_mem_axi_0_b_ready,
  input   io_mem_axi_0_b_valid,
  input  [1:0] io_mem_axi_0_b_bits_resp,
  input  [4:0] io_mem_axi_0_b_bits_id,
  input   io_mem_axi_0_b_bits_user,
  input   io_mem_axi_0_ar_ready,
  output  io_mem_axi_0_ar_valid,
  output [31:0] io_mem_axi_0_ar_bits_addr,
  output [7:0] io_mem_axi_0_ar_bits_len,
  output [2:0] io_mem_axi_0_ar_bits_size,
  output [1:0] io_mem_axi_0_ar_bits_burst,
  output  io_mem_axi_0_ar_bits_lock,
  output [3:0] io_mem_axi_0_ar_bits_cache,
  output [2:0] io_mem_axi_0_ar_bits_prot,
  output [3:0] io_mem_axi_0_ar_bits_qos,
  output [3:0] io_mem_axi_0_ar_bits_region,
  output [4:0] io_mem_axi_0_ar_bits_id,
  output  io_mem_axi_0_ar_bits_user,
  output  io_mem_axi_0_r_ready,
  input   io_mem_axi_0_r_valid,
  input  [1:0] io_mem_axi_0_r_bits_resp,
  input  [63:0] io_mem_axi_0_r_bits_data,
  input   io_mem_axi_0_r_bits_last,
  input  [4:0] io_mem_axi_0_r_bits_id,
  input   io_mem_axi_0_r_bits_user,
  output  io_tiles_cached_0_acquire_ready,
  input   io_tiles_cached_0_acquire_valid,
  input  [25:0] io_tiles_cached_0_acquire_bits_addr_block,
  input   io_tiles_cached_0_acquire_bits_client_xact_id,
  input  [2:0] io_tiles_cached_0_acquire_bits_addr_beat,
  input   io_tiles_cached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_tiles_cached_0_acquire_bits_a_type,
  input  [11:0] io_tiles_cached_0_acquire_bits_union,
  input  [63:0] io_tiles_cached_0_acquire_bits_data,
  input   io_tiles_cached_0_probe_ready,
  output  io_tiles_cached_0_probe_valid,
  output [25:0] io_tiles_cached_0_probe_bits_addr_block,
  output [1:0] io_tiles_cached_0_probe_bits_p_type,
  output  io_tiles_cached_0_release_ready,
  input   io_tiles_cached_0_release_valid,
  input  [2:0] io_tiles_cached_0_release_bits_addr_beat,
  input  [25:0] io_tiles_cached_0_release_bits_addr_block,
  input   io_tiles_cached_0_release_bits_client_xact_id,
  input   io_tiles_cached_0_release_bits_voluntary,
  input  [2:0] io_tiles_cached_0_release_bits_r_type,
  input  [63:0] io_tiles_cached_0_release_bits_data,
  input   io_tiles_cached_0_grant_ready,
  output  io_tiles_cached_0_grant_valid,
  output [2:0] io_tiles_cached_0_grant_bits_addr_beat,
  output  io_tiles_cached_0_grant_bits_client_xact_id,
  output [1:0] io_tiles_cached_0_grant_bits_manager_xact_id,
  output  io_tiles_cached_0_grant_bits_is_builtin_type,
  output [3:0] io_tiles_cached_0_grant_bits_g_type,
  output [63:0] io_tiles_cached_0_grant_bits_data,
  output  io_tiles_cached_0_grant_bits_manager_id,
  output  io_tiles_cached_0_finish_ready,
  input   io_tiles_cached_0_finish_valid,
  input  [1:0] io_tiles_cached_0_finish_bits_manager_xact_id,
  input   io_tiles_cached_0_finish_bits_manager_id,
  output  io_tiles_uncached_0_acquire_ready,
  input   io_tiles_uncached_0_acquire_valid,
  input  [25:0] io_tiles_uncached_0_acquire_bits_addr_block,
  input   io_tiles_uncached_0_acquire_bits_client_xact_id,
  input  [2:0] io_tiles_uncached_0_acquire_bits_addr_beat,
  input   io_tiles_uncached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_tiles_uncached_0_acquire_bits_a_type,
  input  [11:0] io_tiles_uncached_0_acquire_bits_union,
  input  [63:0] io_tiles_uncached_0_acquire_bits_data,
  input   io_tiles_uncached_0_grant_ready,
  output  io_tiles_uncached_0_grant_valid,
  output [2:0] io_tiles_uncached_0_grant_bits_addr_beat,
  output  io_tiles_uncached_0_grant_bits_client_xact_id,
  output [1:0] io_tiles_uncached_0_grant_bits_manager_xact_id,
  output  io_tiles_uncached_0_grant_bits_is_builtin_type,
  output [3:0] io_tiles_uncached_0_grant_bits_g_type,
  output [63:0] io_tiles_uncached_0_grant_bits_data,
  output  io_prci_0_reset,
  output  io_prci_0_id,
  output  io_prci_0_interrupts_meip,
  output  io_prci_0_interrupts_seip,
  output  io_prci_0_interrupts_debug,
  output  io_prci_0_interrupts_mtip,
  output  io_prci_0_interrupts_msip,
  input   io_mmio_axi_0_aw_ready,
  output  io_mmio_axi_0_aw_valid,
  output [31:0] io_mmio_axi_0_aw_bits_addr,
  output [7:0] io_mmio_axi_0_aw_bits_len,
  output [2:0] io_mmio_axi_0_aw_bits_size,
  output [1:0] io_mmio_axi_0_aw_bits_burst,
  output  io_mmio_axi_0_aw_bits_lock,
  output [3:0] io_mmio_axi_0_aw_bits_cache,
  output [2:0] io_mmio_axi_0_aw_bits_prot,
  output [3:0] io_mmio_axi_0_aw_bits_qos,
  output [3:0] io_mmio_axi_0_aw_bits_region,
  output [4:0] io_mmio_axi_0_aw_bits_id,
  output  io_mmio_axi_0_aw_bits_user,
  input   io_mmio_axi_0_w_ready,
  output  io_mmio_axi_0_w_valid,
  output [63:0] io_mmio_axi_0_w_bits_data,
  output  io_mmio_axi_0_w_bits_last,
  output [4:0] io_mmio_axi_0_w_bits_id,
  output [7:0] io_mmio_axi_0_w_bits_strb,
  output  io_mmio_axi_0_w_bits_user,
  output  io_mmio_axi_0_b_ready,
  input   io_mmio_axi_0_b_valid,
  input  [1:0] io_mmio_axi_0_b_bits_resp,
  input  [4:0] io_mmio_axi_0_b_bits_id,
  input   io_mmio_axi_0_b_bits_user,
  input   io_mmio_axi_0_ar_ready,
  output  io_mmio_axi_0_ar_valid,
  output [31:0] io_mmio_axi_0_ar_bits_addr,
  output [7:0] io_mmio_axi_0_ar_bits_len,
  output [2:0] io_mmio_axi_0_ar_bits_size,
  output [1:0] io_mmio_axi_0_ar_bits_burst,
  output  io_mmio_axi_0_ar_bits_lock,
  output [3:0] io_mmio_axi_0_ar_bits_cache,
  output [2:0] io_mmio_axi_0_ar_bits_prot,
  output [3:0] io_mmio_axi_0_ar_bits_qos,
  output [3:0] io_mmio_axi_0_ar_bits_region,
  output [4:0] io_mmio_axi_0_ar_bits_id,
  output  io_mmio_axi_0_ar_bits_user,
  output  io_mmio_axi_0_r_ready,
  input   io_mmio_axi_0_r_valid,
  input  [1:0] io_mmio_axi_0_r_bits_resp,
  input  [63:0] io_mmio_axi_0_r_bits_data,
  input   io_mmio_axi_0_r_bits_last,
  input  [4:0] io_mmio_axi_0_r_bits_id,
  input   io_mmio_axi_0_r_bits_user,
  input   io_interrupts_0,
  input   io_interrupts_1,
  input   io_interrupts_2,
  input   io_interrupts_3,
  input   io_interrupts_4,
  input   io_interrupts_5,
  input   io_interrupts_6,
  input   io_interrupts_7,
  input   io_interrupts_8,
  input   io_interrupts_9,
  input   io_interrupts_10,
  input   io_interrupts_11,
  input   io_interrupts_12,
  input   io_interrupts_13,
  input   io_interrupts_14,
  input   io_interrupts_15,
  input   io_interrupts_16,
  input   io_interrupts_17,
  input   io_interrupts_18,
  input   io_interrupts_19,
  input   io_interrupts_20,
  input   io_interrupts_21,
  input   io_interrupts_22,
  input   io_interrupts_23,
  input   io_interrupts_24,
  input   io_interrupts_25,
  input   io_interrupts_26,
  input   io_interrupts_27,
  input   io_interrupts_28,
  input   io_interrupts_29,
  input   io_interrupts_30,
  output  io_debugBus_req_ready,
  input   io_debugBus_req_valid,
  input  [4:0] io_debugBus_req_bits_addr,
  input  [1:0] io_debugBus_req_bits_op,
  input  [33:0] io_debugBus_req_bits_data,
  input   io_debugBus_resp_ready,
  output  io_debugBus_resp_valid,
  output [1:0] io_debugBus_resp_bits_resp,
  output [33:0] io_debugBus_resp_bits_data
);
  wire  outmemsys_clk;
  wire  outmemsys_reset;
  wire  outmemsys_io_tiles_cached_0_acquire_ready;
  wire  outmemsys_io_tiles_cached_0_acquire_valid;
  wire [25:0] outmemsys_io_tiles_cached_0_acquire_bits_addr_block;
  wire  outmemsys_io_tiles_cached_0_acquire_bits_client_xact_id;
  wire [2:0] outmemsys_io_tiles_cached_0_acquire_bits_addr_beat;
  wire  outmemsys_io_tiles_cached_0_acquire_bits_is_builtin_type;
  wire [2:0] outmemsys_io_tiles_cached_0_acquire_bits_a_type;
  wire [11:0] outmemsys_io_tiles_cached_0_acquire_bits_union;
  wire [63:0] outmemsys_io_tiles_cached_0_acquire_bits_data;
  wire  outmemsys_io_tiles_cached_0_probe_ready;
  wire  outmemsys_io_tiles_cached_0_probe_valid;
  wire [25:0] outmemsys_io_tiles_cached_0_probe_bits_addr_block;
  wire [1:0] outmemsys_io_tiles_cached_0_probe_bits_p_type;
  wire  outmemsys_io_tiles_cached_0_release_ready;
  wire  outmemsys_io_tiles_cached_0_release_valid;
  wire [2:0] outmemsys_io_tiles_cached_0_release_bits_addr_beat;
  wire [25:0] outmemsys_io_tiles_cached_0_release_bits_addr_block;
  wire  outmemsys_io_tiles_cached_0_release_bits_client_xact_id;
  wire  outmemsys_io_tiles_cached_0_release_bits_voluntary;
  wire [2:0] outmemsys_io_tiles_cached_0_release_bits_r_type;
  wire [63:0] outmemsys_io_tiles_cached_0_release_bits_data;
  wire  outmemsys_io_tiles_cached_0_grant_ready;
  wire  outmemsys_io_tiles_cached_0_grant_valid;
  wire [2:0] outmemsys_io_tiles_cached_0_grant_bits_addr_beat;
  wire  outmemsys_io_tiles_cached_0_grant_bits_client_xact_id;
  wire [1:0] outmemsys_io_tiles_cached_0_grant_bits_manager_xact_id;
  wire  outmemsys_io_tiles_cached_0_grant_bits_is_builtin_type;
  wire [3:0] outmemsys_io_tiles_cached_0_grant_bits_g_type;
  wire [63:0] outmemsys_io_tiles_cached_0_grant_bits_data;
  wire  outmemsys_io_tiles_cached_0_grant_bits_manager_id;
  wire  outmemsys_io_tiles_cached_0_finish_ready;
  wire  outmemsys_io_tiles_cached_0_finish_valid;
  wire [1:0] outmemsys_io_tiles_cached_0_finish_bits_manager_xact_id;
  wire  outmemsys_io_tiles_cached_0_finish_bits_manager_id;
  wire  outmemsys_io_tiles_uncached_0_acquire_ready;
  wire  outmemsys_io_tiles_uncached_0_acquire_valid;
  wire [25:0] outmemsys_io_tiles_uncached_0_acquire_bits_addr_block;
  wire  outmemsys_io_tiles_uncached_0_acquire_bits_client_xact_id;
  wire [2:0] outmemsys_io_tiles_uncached_0_acquire_bits_addr_beat;
  wire  outmemsys_io_tiles_uncached_0_acquire_bits_is_builtin_type;
  wire [2:0] outmemsys_io_tiles_uncached_0_acquire_bits_a_type;
  wire [11:0] outmemsys_io_tiles_uncached_0_acquire_bits_union;
  wire [63:0] outmemsys_io_tiles_uncached_0_acquire_bits_data;
  wire  outmemsys_io_tiles_uncached_0_grant_ready;
  wire  outmemsys_io_tiles_uncached_0_grant_valid;
  wire [2:0] outmemsys_io_tiles_uncached_0_grant_bits_addr_beat;
  wire  outmemsys_io_tiles_uncached_0_grant_bits_client_xact_id;
  wire [1:0] outmemsys_io_tiles_uncached_0_grant_bits_manager_xact_id;
  wire  outmemsys_io_tiles_uncached_0_grant_bits_is_builtin_type;
  wire [3:0] outmemsys_io_tiles_uncached_0_grant_bits_g_type;
  wire [63:0] outmemsys_io_tiles_uncached_0_grant_bits_data;
  wire  outmemsys_io_incoherent_0;
  wire  outmemsys_io_mem_axi_0_aw_ready;
  wire  outmemsys_io_mem_axi_0_aw_valid;
  wire [31:0] outmemsys_io_mem_axi_0_aw_bits_addr;
  wire [7:0] outmemsys_io_mem_axi_0_aw_bits_len;
  wire [2:0] outmemsys_io_mem_axi_0_aw_bits_size;
  wire [1:0] outmemsys_io_mem_axi_0_aw_bits_burst;
  wire  outmemsys_io_mem_axi_0_aw_bits_lock;
  wire [3:0] outmemsys_io_mem_axi_0_aw_bits_cache;
  wire [2:0] outmemsys_io_mem_axi_0_aw_bits_prot;
  wire [3:0] outmemsys_io_mem_axi_0_aw_bits_qos;
  wire [3:0] outmemsys_io_mem_axi_0_aw_bits_region;
  wire [4:0] outmemsys_io_mem_axi_0_aw_bits_id;
  wire  outmemsys_io_mem_axi_0_aw_bits_user;
  wire  outmemsys_io_mem_axi_0_w_ready;
  wire  outmemsys_io_mem_axi_0_w_valid;
  wire [63:0] outmemsys_io_mem_axi_0_w_bits_data;
  wire  outmemsys_io_mem_axi_0_w_bits_last;
  wire [4:0] outmemsys_io_mem_axi_0_w_bits_id;
  wire [7:0] outmemsys_io_mem_axi_0_w_bits_strb;
  wire  outmemsys_io_mem_axi_0_w_bits_user;
  wire  outmemsys_io_mem_axi_0_b_ready;
  wire  outmemsys_io_mem_axi_0_b_valid;
  wire [1:0] outmemsys_io_mem_axi_0_b_bits_resp;
  wire [4:0] outmemsys_io_mem_axi_0_b_bits_id;
  wire  outmemsys_io_mem_axi_0_b_bits_user;
  wire  outmemsys_io_mem_axi_0_ar_ready;
  wire  outmemsys_io_mem_axi_0_ar_valid;
  wire [31:0] outmemsys_io_mem_axi_0_ar_bits_addr;
  wire [7:0] outmemsys_io_mem_axi_0_ar_bits_len;
  wire [2:0] outmemsys_io_mem_axi_0_ar_bits_size;
  wire [1:0] outmemsys_io_mem_axi_0_ar_bits_burst;
  wire  outmemsys_io_mem_axi_0_ar_bits_lock;
  wire [3:0] outmemsys_io_mem_axi_0_ar_bits_cache;
  wire [2:0] outmemsys_io_mem_axi_0_ar_bits_prot;
  wire [3:0] outmemsys_io_mem_axi_0_ar_bits_qos;
  wire [3:0] outmemsys_io_mem_axi_0_ar_bits_region;
  wire [4:0] outmemsys_io_mem_axi_0_ar_bits_id;
  wire  outmemsys_io_mem_axi_0_ar_bits_user;
  wire  outmemsys_io_mem_axi_0_r_ready;
  wire  outmemsys_io_mem_axi_0_r_valid;
  wire [1:0] outmemsys_io_mem_axi_0_r_bits_resp;
  wire [63:0] outmemsys_io_mem_axi_0_r_bits_data;
  wire  outmemsys_io_mem_axi_0_r_bits_last;
  wire [4:0] outmemsys_io_mem_axi_0_r_bits_id;
  wire  outmemsys_io_mem_axi_0_r_bits_user;
  wire  outmemsys_io_mmio_acquire_ready;
  wire  outmemsys_io_mmio_acquire_valid;
  wire [25:0] outmemsys_io_mmio_acquire_bits_addr_block;
  wire [1:0] outmemsys_io_mmio_acquire_bits_client_xact_id;
  wire [2:0] outmemsys_io_mmio_acquire_bits_addr_beat;
  wire  outmemsys_io_mmio_acquire_bits_is_builtin_type;
  wire [2:0] outmemsys_io_mmio_acquire_bits_a_type;
  wire [11:0] outmemsys_io_mmio_acquire_bits_union;
  wire [63:0] outmemsys_io_mmio_acquire_bits_data;
  wire  outmemsys_io_mmio_grant_ready;
  wire  outmemsys_io_mmio_grant_valid;
  wire [2:0] outmemsys_io_mmio_grant_bits_addr_beat;
  wire [1:0] outmemsys_io_mmio_grant_bits_client_xact_id;
  wire  outmemsys_io_mmio_grant_bits_manager_xact_id;
  wire  outmemsys_io_mmio_grant_bits_is_builtin_type;
  wire [3:0] outmemsys_io_mmio_grant_bits_g_type;
  wire [63:0] outmemsys_io_mmio_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_clk;
  wire  TileLinkRecursiveInterconnect_2_reset;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_4_acquire_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_4_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_2_io_out_4_grant_ready;
  wire  TileLinkRecursiveInterconnect_2_io_out_4_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_data;
  wire  PLIC_1_clk;
  wire  PLIC_1_reset;
  wire  PLIC_1_io_devices_0_valid;
  wire  PLIC_1_io_devices_0_ready;
  wire  PLIC_1_io_devices_0_complete;
  wire  PLIC_1_io_devices_1_valid;
  wire  PLIC_1_io_devices_1_ready;
  wire  PLIC_1_io_devices_1_complete;
  wire  PLIC_1_io_devices_2_valid;
  wire  PLIC_1_io_devices_2_ready;
  wire  PLIC_1_io_devices_2_complete;
  wire  PLIC_1_io_devices_3_valid;
  wire  PLIC_1_io_devices_3_ready;
  wire  PLIC_1_io_devices_3_complete;
  wire  PLIC_1_io_devices_4_valid;
  wire  PLIC_1_io_devices_4_ready;
  wire  PLIC_1_io_devices_4_complete;
  wire  PLIC_1_io_devices_5_valid;
  wire  PLIC_1_io_devices_5_ready;
  wire  PLIC_1_io_devices_5_complete;
  wire  PLIC_1_io_devices_6_valid;
  wire  PLIC_1_io_devices_6_ready;
  wire  PLIC_1_io_devices_6_complete;
  wire  PLIC_1_io_devices_7_valid;
  wire  PLIC_1_io_devices_7_ready;
  wire  PLIC_1_io_devices_7_complete;
  wire  PLIC_1_io_devices_8_valid;
  wire  PLIC_1_io_devices_8_ready;
  wire  PLIC_1_io_devices_8_complete;
  wire  PLIC_1_io_devices_9_valid;
  wire  PLIC_1_io_devices_9_ready;
  wire  PLIC_1_io_devices_9_complete;
  wire  PLIC_1_io_devices_10_valid;
  wire  PLIC_1_io_devices_10_ready;
  wire  PLIC_1_io_devices_10_complete;
  wire  PLIC_1_io_devices_11_valid;
  wire  PLIC_1_io_devices_11_ready;
  wire  PLIC_1_io_devices_11_complete;
  wire  PLIC_1_io_devices_12_valid;
  wire  PLIC_1_io_devices_12_ready;
  wire  PLIC_1_io_devices_12_complete;
  wire  PLIC_1_io_devices_13_valid;
  wire  PLIC_1_io_devices_13_ready;
  wire  PLIC_1_io_devices_13_complete;
  wire  PLIC_1_io_devices_14_valid;
  wire  PLIC_1_io_devices_14_ready;
  wire  PLIC_1_io_devices_14_complete;
  wire  PLIC_1_io_devices_15_valid;
  wire  PLIC_1_io_devices_15_ready;
  wire  PLIC_1_io_devices_15_complete;
  wire  PLIC_1_io_devices_16_valid;
  wire  PLIC_1_io_devices_16_ready;
  wire  PLIC_1_io_devices_16_complete;
  wire  PLIC_1_io_devices_17_valid;
  wire  PLIC_1_io_devices_17_ready;
  wire  PLIC_1_io_devices_17_complete;
  wire  PLIC_1_io_devices_18_valid;
  wire  PLIC_1_io_devices_18_ready;
  wire  PLIC_1_io_devices_18_complete;
  wire  PLIC_1_io_devices_19_valid;
  wire  PLIC_1_io_devices_19_ready;
  wire  PLIC_1_io_devices_19_complete;
  wire  PLIC_1_io_devices_20_valid;
  wire  PLIC_1_io_devices_20_ready;
  wire  PLIC_1_io_devices_20_complete;
  wire  PLIC_1_io_devices_21_valid;
  wire  PLIC_1_io_devices_21_ready;
  wire  PLIC_1_io_devices_21_complete;
  wire  PLIC_1_io_devices_22_valid;
  wire  PLIC_1_io_devices_22_ready;
  wire  PLIC_1_io_devices_22_complete;
  wire  PLIC_1_io_devices_23_valid;
  wire  PLIC_1_io_devices_23_ready;
  wire  PLIC_1_io_devices_23_complete;
  wire  PLIC_1_io_devices_24_valid;
  wire  PLIC_1_io_devices_24_ready;
  wire  PLIC_1_io_devices_24_complete;
  wire  PLIC_1_io_devices_25_valid;
  wire  PLIC_1_io_devices_25_ready;
  wire  PLIC_1_io_devices_25_complete;
  wire  PLIC_1_io_devices_26_valid;
  wire  PLIC_1_io_devices_26_ready;
  wire  PLIC_1_io_devices_26_complete;
  wire  PLIC_1_io_devices_27_valid;
  wire  PLIC_1_io_devices_27_ready;
  wire  PLIC_1_io_devices_27_complete;
  wire  PLIC_1_io_devices_28_valid;
  wire  PLIC_1_io_devices_28_ready;
  wire  PLIC_1_io_devices_28_complete;
  wire  PLIC_1_io_devices_29_valid;
  wire  PLIC_1_io_devices_29_ready;
  wire  PLIC_1_io_devices_29_complete;
  wire  PLIC_1_io_devices_30_valid;
  wire  PLIC_1_io_devices_30_ready;
  wire  PLIC_1_io_devices_30_complete;
  wire  PLIC_1_io_harts_0;
  wire  PLIC_1_io_tl_acquire_ready;
  wire  PLIC_1_io_tl_acquire_valid;
  wire [25:0] PLIC_1_io_tl_acquire_bits_addr_block;
  wire [1:0] PLIC_1_io_tl_acquire_bits_client_xact_id;
  wire [2:0] PLIC_1_io_tl_acquire_bits_addr_beat;
  wire  PLIC_1_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] PLIC_1_io_tl_acquire_bits_a_type;
  wire [11:0] PLIC_1_io_tl_acquire_bits_union;
  wire [63:0] PLIC_1_io_tl_acquire_bits_data;
  wire  PLIC_1_io_tl_grant_ready;
  wire  PLIC_1_io_tl_grant_valid;
  wire [2:0] PLIC_1_io_tl_grant_bits_addr_beat;
  wire [1:0] PLIC_1_io_tl_grant_bits_client_xact_id;
  wire  PLIC_1_io_tl_grant_bits_manager_xact_id;
  wire  PLIC_1_io_tl_grant_bits_is_builtin_type;
  wire [3:0] PLIC_1_io_tl_grant_bits_g_type;
  wire [63:0] PLIC_1_io_tl_grant_bits_data;
  wire  LevelGateway_31_clk;
  wire  LevelGateway_31_reset;
  wire  LevelGateway_31_io_interrupt;
  wire  LevelGateway_31_io_plic_valid;
  wire  LevelGateway_31_io_plic_ready;
  wire  LevelGateway_31_io_plic_complete;
  wire  LevelGateway_1_1_clk;
  wire  LevelGateway_1_1_reset;
  wire  LevelGateway_1_1_io_interrupt;
  wire  LevelGateway_1_1_io_plic_valid;
  wire  LevelGateway_1_1_io_plic_ready;
  wire  LevelGateway_1_1_io_plic_complete;
  wire  LevelGateway_2_1_clk;
  wire  LevelGateway_2_1_reset;
  wire  LevelGateway_2_1_io_interrupt;
  wire  LevelGateway_2_1_io_plic_valid;
  wire  LevelGateway_2_1_io_plic_ready;
  wire  LevelGateway_2_1_io_plic_complete;
  wire  LevelGateway_3_1_clk;
  wire  LevelGateway_3_1_reset;
  wire  LevelGateway_3_1_io_interrupt;
  wire  LevelGateway_3_1_io_plic_valid;
  wire  LevelGateway_3_1_io_plic_ready;
  wire  LevelGateway_3_1_io_plic_complete;
  wire  LevelGateway_4_1_clk;
  wire  LevelGateway_4_1_reset;
  wire  LevelGateway_4_1_io_interrupt;
  wire  LevelGateway_4_1_io_plic_valid;
  wire  LevelGateway_4_1_io_plic_ready;
  wire  LevelGateway_4_1_io_plic_complete;
  wire  LevelGateway_5_1_clk;
  wire  LevelGateway_5_1_reset;
  wire  LevelGateway_5_1_io_interrupt;
  wire  LevelGateway_5_1_io_plic_valid;
  wire  LevelGateway_5_1_io_plic_ready;
  wire  LevelGateway_5_1_io_plic_complete;
  wire  LevelGateway_6_1_clk;
  wire  LevelGateway_6_1_reset;
  wire  LevelGateway_6_1_io_interrupt;
  wire  LevelGateway_6_1_io_plic_valid;
  wire  LevelGateway_6_1_io_plic_ready;
  wire  LevelGateway_6_1_io_plic_complete;
  wire  LevelGateway_7_1_clk;
  wire  LevelGateway_7_1_reset;
  wire  LevelGateway_7_1_io_interrupt;
  wire  LevelGateway_7_1_io_plic_valid;
  wire  LevelGateway_7_1_io_plic_ready;
  wire  LevelGateway_7_1_io_plic_complete;
  wire  LevelGateway_8_1_clk;
  wire  LevelGateway_8_1_reset;
  wire  LevelGateway_8_1_io_interrupt;
  wire  LevelGateway_8_1_io_plic_valid;
  wire  LevelGateway_8_1_io_plic_ready;
  wire  LevelGateway_8_1_io_plic_complete;
  wire  LevelGateway_9_1_clk;
  wire  LevelGateway_9_1_reset;
  wire  LevelGateway_9_1_io_interrupt;
  wire  LevelGateway_9_1_io_plic_valid;
  wire  LevelGateway_9_1_io_plic_ready;
  wire  LevelGateway_9_1_io_plic_complete;
  wire  LevelGateway_10_1_clk;
  wire  LevelGateway_10_1_reset;
  wire  LevelGateway_10_1_io_interrupt;
  wire  LevelGateway_10_1_io_plic_valid;
  wire  LevelGateway_10_1_io_plic_ready;
  wire  LevelGateway_10_1_io_plic_complete;
  wire  LevelGateway_11_1_clk;
  wire  LevelGateway_11_1_reset;
  wire  LevelGateway_11_1_io_interrupt;
  wire  LevelGateway_11_1_io_plic_valid;
  wire  LevelGateway_11_1_io_plic_ready;
  wire  LevelGateway_11_1_io_plic_complete;
  wire  LevelGateway_12_1_clk;
  wire  LevelGateway_12_1_reset;
  wire  LevelGateway_12_1_io_interrupt;
  wire  LevelGateway_12_1_io_plic_valid;
  wire  LevelGateway_12_1_io_plic_ready;
  wire  LevelGateway_12_1_io_plic_complete;
  wire  LevelGateway_13_1_clk;
  wire  LevelGateway_13_1_reset;
  wire  LevelGateway_13_1_io_interrupt;
  wire  LevelGateway_13_1_io_plic_valid;
  wire  LevelGateway_13_1_io_plic_ready;
  wire  LevelGateway_13_1_io_plic_complete;
  wire  LevelGateway_14_1_clk;
  wire  LevelGateway_14_1_reset;
  wire  LevelGateway_14_1_io_interrupt;
  wire  LevelGateway_14_1_io_plic_valid;
  wire  LevelGateway_14_1_io_plic_ready;
  wire  LevelGateway_14_1_io_plic_complete;
  wire  LevelGateway_15_1_clk;
  wire  LevelGateway_15_1_reset;
  wire  LevelGateway_15_1_io_interrupt;
  wire  LevelGateway_15_1_io_plic_valid;
  wire  LevelGateway_15_1_io_plic_ready;
  wire  LevelGateway_15_1_io_plic_complete;
  wire  LevelGateway_16_1_clk;
  wire  LevelGateway_16_1_reset;
  wire  LevelGateway_16_1_io_interrupt;
  wire  LevelGateway_16_1_io_plic_valid;
  wire  LevelGateway_16_1_io_plic_ready;
  wire  LevelGateway_16_1_io_plic_complete;
  wire  LevelGateway_17_1_clk;
  wire  LevelGateway_17_1_reset;
  wire  LevelGateway_17_1_io_interrupt;
  wire  LevelGateway_17_1_io_plic_valid;
  wire  LevelGateway_17_1_io_plic_ready;
  wire  LevelGateway_17_1_io_plic_complete;
  wire  LevelGateway_18_1_clk;
  wire  LevelGateway_18_1_reset;
  wire  LevelGateway_18_1_io_interrupt;
  wire  LevelGateway_18_1_io_plic_valid;
  wire  LevelGateway_18_1_io_plic_ready;
  wire  LevelGateway_18_1_io_plic_complete;
  wire  LevelGateway_19_1_clk;
  wire  LevelGateway_19_1_reset;
  wire  LevelGateway_19_1_io_interrupt;
  wire  LevelGateway_19_1_io_plic_valid;
  wire  LevelGateway_19_1_io_plic_ready;
  wire  LevelGateway_19_1_io_plic_complete;
  wire  LevelGateway_20_1_clk;
  wire  LevelGateway_20_1_reset;
  wire  LevelGateway_20_1_io_interrupt;
  wire  LevelGateway_20_1_io_plic_valid;
  wire  LevelGateway_20_1_io_plic_ready;
  wire  LevelGateway_20_1_io_plic_complete;
  wire  LevelGateway_21_1_clk;
  wire  LevelGateway_21_1_reset;
  wire  LevelGateway_21_1_io_interrupt;
  wire  LevelGateway_21_1_io_plic_valid;
  wire  LevelGateway_21_1_io_plic_ready;
  wire  LevelGateway_21_1_io_plic_complete;
  wire  LevelGateway_22_1_clk;
  wire  LevelGateway_22_1_reset;
  wire  LevelGateway_22_1_io_interrupt;
  wire  LevelGateway_22_1_io_plic_valid;
  wire  LevelGateway_22_1_io_plic_ready;
  wire  LevelGateway_22_1_io_plic_complete;
  wire  LevelGateway_23_1_clk;
  wire  LevelGateway_23_1_reset;
  wire  LevelGateway_23_1_io_interrupt;
  wire  LevelGateway_23_1_io_plic_valid;
  wire  LevelGateway_23_1_io_plic_ready;
  wire  LevelGateway_23_1_io_plic_complete;
  wire  LevelGateway_24_1_clk;
  wire  LevelGateway_24_1_reset;
  wire  LevelGateway_24_1_io_interrupt;
  wire  LevelGateway_24_1_io_plic_valid;
  wire  LevelGateway_24_1_io_plic_ready;
  wire  LevelGateway_24_1_io_plic_complete;
  wire  LevelGateway_25_1_clk;
  wire  LevelGateway_25_1_reset;
  wire  LevelGateway_25_1_io_interrupt;
  wire  LevelGateway_25_1_io_plic_valid;
  wire  LevelGateway_25_1_io_plic_ready;
  wire  LevelGateway_25_1_io_plic_complete;
  wire  LevelGateway_26_1_clk;
  wire  LevelGateway_26_1_reset;
  wire  LevelGateway_26_1_io_interrupt;
  wire  LevelGateway_26_1_io_plic_valid;
  wire  LevelGateway_26_1_io_plic_ready;
  wire  LevelGateway_26_1_io_plic_complete;
  wire  LevelGateway_27_1_clk;
  wire  LevelGateway_27_1_reset;
  wire  LevelGateway_27_1_io_interrupt;
  wire  LevelGateway_27_1_io_plic_valid;
  wire  LevelGateway_27_1_io_plic_ready;
  wire  LevelGateway_27_1_io_plic_complete;
  wire  LevelGateway_28_1_clk;
  wire  LevelGateway_28_1_reset;
  wire  LevelGateway_28_1_io_interrupt;
  wire  LevelGateway_28_1_io_plic_valid;
  wire  LevelGateway_28_1_io_plic_ready;
  wire  LevelGateway_28_1_io_plic_complete;
  wire  LevelGateway_29_1_clk;
  wire  LevelGateway_29_1_reset;
  wire  LevelGateway_29_1_io_interrupt;
  wire  LevelGateway_29_1_io_plic_valid;
  wire  LevelGateway_29_1_io_plic_ready;
  wire  LevelGateway_29_1_io_plic_complete;
  wire  LevelGateway_30_1_clk;
  wire  LevelGateway_30_1_reset;
  wire  LevelGateway_30_1_io_interrupt;
  wire  LevelGateway_30_1_io_plic_valid;
  wire  LevelGateway_30_1_io_plic_ready;
  wire  LevelGateway_30_1_io_plic_complete;
  wire  DebugModule_1_clk;
  wire  DebugModule_1_reset;
  wire  DebugModule_1_io_db_req_ready;
  wire  DebugModule_1_io_db_req_valid;
  wire [4:0] DebugModule_1_io_db_req_bits_addr;
  wire [1:0] DebugModule_1_io_db_req_bits_op;
  wire [33:0] DebugModule_1_io_db_req_bits_data;
  wire  DebugModule_1_io_db_resp_ready;
  wire  DebugModule_1_io_db_resp_valid;
  wire [1:0] DebugModule_1_io_db_resp_bits_resp;
  wire [33:0] DebugModule_1_io_db_resp_bits_data;
  wire  DebugModule_1_io_debugInterrupts_0;
  wire  DebugModule_1_io_tl_acquire_ready;
  wire  DebugModule_1_io_tl_acquire_valid;
  wire [25:0] DebugModule_1_io_tl_acquire_bits_addr_block;
  wire [1:0] DebugModule_1_io_tl_acquire_bits_client_xact_id;
  wire [2:0] DebugModule_1_io_tl_acquire_bits_addr_beat;
  wire  DebugModule_1_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] DebugModule_1_io_tl_acquire_bits_a_type;
  wire [11:0] DebugModule_1_io_tl_acquire_bits_union;
  wire [63:0] DebugModule_1_io_tl_acquire_bits_data;
  wire  DebugModule_1_io_tl_grant_ready;
  wire  DebugModule_1_io_tl_grant_valid;
  wire [2:0] DebugModule_1_io_tl_grant_bits_addr_beat;
  wire [1:0] DebugModule_1_io_tl_grant_bits_client_xact_id;
  wire  DebugModule_1_io_tl_grant_bits_manager_xact_id;
  wire  DebugModule_1_io_tl_grant_bits_is_builtin_type;
  wire [3:0] DebugModule_1_io_tl_grant_bits_g_type;
  wire [63:0] DebugModule_1_io_tl_grant_bits_data;
  wire  DebugModule_1_io_ndreset;
  wire  DebugModule_1_io_fullreset;
  wire  PRCI_1_clk;
  wire  PRCI_1_reset;
  wire  PRCI_1_io_interrupts_0_meip;
  wire  PRCI_1_io_interrupts_0_seip;
  wire  PRCI_1_io_interrupts_0_debug;
  wire  PRCI_1_io_tl_acquire_ready;
  wire  PRCI_1_io_tl_acquire_valid;
  wire [25:0] PRCI_1_io_tl_acquire_bits_addr_block;
  wire [1:0] PRCI_1_io_tl_acquire_bits_client_xact_id;
  wire [2:0] PRCI_1_io_tl_acquire_bits_addr_beat;
  wire  PRCI_1_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] PRCI_1_io_tl_acquire_bits_a_type;
  wire [11:0] PRCI_1_io_tl_acquire_bits_union;
  wire [63:0] PRCI_1_io_tl_acquire_bits_data;
  wire  PRCI_1_io_tl_grant_ready;
  wire  PRCI_1_io_tl_grant_valid;
  wire [2:0] PRCI_1_io_tl_grant_bits_addr_beat;
  wire [1:0] PRCI_1_io_tl_grant_bits_client_xact_id;
  wire  PRCI_1_io_tl_grant_bits_manager_xact_id;
  wire  PRCI_1_io_tl_grant_bits_is_builtin_type;
  wire [3:0] PRCI_1_io_tl_grant_bits_g_type;
  wire [63:0] PRCI_1_io_tl_grant_bits_data;
  wire  PRCI_1_io_tiles_0_reset;
  wire  PRCI_1_io_tiles_0_id;
  wire  PRCI_1_io_tiles_0_interrupts_meip;
  wire  PRCI_1_io_tiles_0_interrupts_seip;
  wire  PRCI_1_io_tiles_0_interrupts_debug;
  wire  PRCI_1_io_tiles_0_interrupts_mtip;
  wire  PRCI_1_io_tiles_0_interrupts_msip;
  wire  PRCI_1_io_rtcTick;
  reg [6:0] T_10389;
  reg [31:0] GEN_2;
  wire  T_10391;
  wire [7:0] T_10393;
  wire [6:0] T_10394;
  wire [6:0] GEN_0;
  wire  ROMSlave_1_clk;
  wire  ROMSlave_1_reset;
  wire  ROMSlave_1_io_acquire_ready;
  wire  ROMSlave_1_io_acquire_valid;
  wire [25:0] ROMSlave_1_io_acquire_bits_addr_block;
  wire [1:0] ROMSlave_1_io_acquire_bits_client_xact_id;
  wire [2:0] ROMSlave_1_io_acquire_bits_addr_beat;
  wire  ROMSlave_1_io_acquire_bits_is_builtin_type;
  wire [2:0] ROMSlave_1_io_acquire_bits_a_type;
  wire [11:0] ROMSlave_1_io_acquire_bits_union;
  wire [63:0] ROMSlave_1_io_acquire_bits_data;
  wire  ROMSlave_1_io_grant_ready;
  wire  ROMSlave_1_io_grant_valid;
  wire [2:0] ROMSlave_1_io_grant_bits_addr_beat;
  wire [1:0] ROMSlave_1_io_grant_bits_client_xact_id;
  wire  ROMSlave_1_io_grant_bits_manager_xact_id;
  wire  ROMSlave_1_io_grant_bits_is_builtin_type;
  wire [3:0] ROMSlave_1_io_grant_bits_g_type;
  wire [63:0] ROMSlave_1_io_grant_bits_data;
  wire  NastiIOTileLinkIOConverter_1_1_clk;
  wire  NastiIOTileLinkIOConverter_1_1_reset;
  wire  NastiIOTileLinkIOConverter_1_1_io_tl_acquire_ready;
  wire  NastiIOTileLinkIOConverter_1_1_io_tl_acquire_valid;
  wire [25:0] NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_addr_block;
  wire [1:0] NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_client_xact_id;
  wire [2:0] NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_addr_beat;
  wire  NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_a_type;
  wire [11:0] NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_union;
  wire [63:0] NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_data;
  wire  NastiIOTileLinkIOConverter_1_1_io_tl_grant_ready;
  wire  NastiIOTileLinkIOConverter_1_1_io_tl_grant_valid;
  wire [2:0] NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_addr_beat;
  wire [1:0] NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_client_xact_id;
  wire  NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_manager_xact_id;
  wire  NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_is_builtin_type;
  wire [3:0] NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_g_type;
  wire [63:0] NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_data;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_aw_ready;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_aw_valid;
  wire [31:0] NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_addr;
  wire [7:0] NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_len;
  wire [2:0] NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_size;
  wire [1:0] NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_burst;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_lock;
  wire [3:0] NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_cache;
  wire [2:0] NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_prot;
  wire [3:0] NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_qos;
  wire [3:0] NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_region;
  wire [4:0] NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_id;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_user;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_w_ready;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_w_valid;
  wire [63:0] NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_data;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_last;
  wire [4:0] NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_id;
  wire [7:0] NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_strb;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_user;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_b_ready;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_b_valid;
  wire [1:0] NastiIOTileLinkIOConverter_1_1_io_nasti_b_bits_resp;
  wire [4:0] NastiIOTileLinkIOConverter_1_1_io_nasti_b_bits_id;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_b_bits_user;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_ar_ready;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_ar_valid;
  wire [31:0] NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_addr;
  wire [7:0] NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_len;
  wire [2:0] NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_size;
  wire [1:0] NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_burst;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_lock;
  wire [3:0] NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_cache;
  wire [2:0] NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_prot;
  wire [3:0] NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_qos;
  wire [3:0] NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_region;
  wire [4:0] NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_id;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_user;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_r_ready;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_r_valid;
  wire [1:0] NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_resp;
  wire [63:0] NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_data;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_last;
  wire [4:0] NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_id;
  wire  NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_user;
  wire  Queue_18_1_clk;
  wire  Queue_18_1_reset;
  wire  Queue_18_1_io_enq_ready;
  wire  Queue_18_1_io_enq_valid;
  wire [31:0] Queue_18_1_io_enq_bits_addr;
  wire [7:0] Queue_18_1_io_enq_bits_len;
  wire [2:0] Queue_18_1_io_enq_bits_size;
  wire [1:0] Queue_18_1_io_enq_bits_burst;
  wire  Queue_18_1_io_enq_bits_lock;
  wire [3:0] Queue_18_1_io_enq_bits_cache;
  wire [2:0] Queue_18_1_io_enq_bits_prot;
  wire [3:0] Queue_18_1_io_enq_bits_qos;
  wire [3:0] Queue_18_1_io_enq_bits_region;
  wire [4:0] Queue_18_1_io_enq_bits_id;
  wire  Queue_18_1_io_enq_bits_user;
  wire  Queue_18_1_io_deq_ready;
  wire  Queue_18_1_io_deq_valid;
  wire [31:0] Queue_18_1_io_deq_bits_addr;
  wire [7:0] Queue_18_1_io_deq_bits_len;
  wire [2:0] Queue_18_1_io_deq_bits_size;
  wire [1:0] Queue_18_1_io_deq_bits_burst;
  wire  Queue_18_1_io_deq_bits_lock;
  wire [3:0] Queue_18_1_io_deq_bits_cache;
  wire [2:0] Queue_18_1_io_deq_bits_prot;
  wire [3:0] Queue_18_1_io_deq_bits_qos;
  wire [3:0] Queue_18_1_io_deq_bits_region;
  wire [4:0] Queue_18_1_io_deq_bits_id;
  wire  Queue_18_1_io_deq_bits_user;
  wire  Queue_18_1_io_count;
  wire  Queue_19_1_clk;
  wire  Queue_19_1_reset;
  wire  Queue_19_1_io_enq_ready;
  wire  Queue_19_1_io_enq_valid;
  wire [31:0] Queue_19_1_io_enq_bits_addr;
  wire [7:0] Queue_19_1_io_enq_bits_len;
  wire [2:0] Queue_19_1_io_enq_bits_size;
  wire [1:0] Queue_19_1_io_enq_bits_burst;
  wire  Queue_19_1_io_enq_bits_lock;
  wire [3:0] Queue_19_1_io_enq_bits_cache;
  wire [2:0] Queue_19_1_io_enq_bits_prot;
  wire [3:0] Queue_19_1_io_enq_bits_qos;
  wire [3:0] Queue_19_1_io_enq_bits_region;
  wire [4:0] Queue_19_1_io_enq_bits_id;
  wire  Queue_19_1_io_enq_bits_user;
  wire  Queue_19_1_io_deq_ready;
  wire  Queue_19_1_io_deq_valid;
  wire [31:0] Queue_19_1_io_deq_bits_addr;
  wire [7:0] Queue_19_1_io_deq_bits_len;
  wire [2:0] Queue_19_1_io_deq_bits_size;
  wire [1:0] Queue_19_1_io_deq_bits_burst;
  wire  Queue_19_1_io_deq_bits_lock;
  wire [3:0] Queue_19_1_io_deq_bits_cache;
  wire [2:0] Queue_19_1_io_deq_bits_prot;
  wire [3:0] Queue_19_1_io_deq_bits_qos;
  wire [3:0] Queue_19_1_io_deq_bits_region;
  wire [4:0] Queue_19_1_io_deq_bits_id;
  wire  Queue_19_1_io_deq_bits_user;
  wire  Queue_19_1_io_count;
  wire  Queue_20_1_clk;
  wire  Queue_20_1_reset;
  wire  Queue_20_1_io_enq_ready;
  wire  Queue_20_1_io_enq_valid;
  wire [63:0] Queue_20_1_io_enq_bits_data;
  wire  Queue_20_1_io_enq_bits_last;
  wire [4:0] Queue_20_1_io_enq_bits_id;
  wire [7:0] Queue_20_1_io_enq_bits_strb;
  wire  Queue_20_1_io_enq_bits_user;
  wire  Queue_20_1_io_deq_ready;
  wire  Queue_20_1_io_deq_valid;
  wire [63:0] Queue_20_1_io_deq_bits_data;
  wire  Queue_20_1_io_deq_bits_last;
  wire [4:0] Queue_20_1_io_deq_bits_id;
  wire [7:0] Queue_20_1_io_deq_bits_strb;
  wire  Queue_20_1_io_deq_bits_user;
  wire [1:0] Queue_20_1_io_count;
  wire  Queue_21_1_clk;
  wire  Queue_21_1_reset;
  wire  Queue_21_1_io_enq_ready;
  wire  Queue_21_1_io_enq_valid;
  wire [1:0] Queue_21_1_io_enq_bits_resp;
  wire [63:0] Queue_21_1_io_enq_bits_data;
  wire  Queue_21_1_io_enq_bits_last;
  wire [4:0] Queue_21_1_io_enq_bits_id;
  wire  Queue_21_1_io_enq_bits_user;
  wire  Queue_21_1_io_deq_ready;
  wire  Queue_21_1_io_deq_valid;
  wire [1:0] Queue_21_1_io_deq_bits_resp;
  wire [63:0] Queue_21_1_io_deq_bits_data;
  wire  Queue_21_1_io_deq_bits_last;
  wire [4:0] Queue_21_1_io_deq_bits_id;
  wire  Queue_21_1_io_deq_bits_user;
  wire [1:0] Queue_21_1_io_count;
  wire  Queue_22_1_clk;
  wire  Queue_22_1_reset;
  wire  Queue_22_1_io_enq_ready;
  wire  Queue_22_1_io_enq_valid;
  wire [1:0] Queue_22_1_io_enq_bits_resp;
  wire [4:0] Queue_22_1_io_enq_bits_id;
  wire  Queue_22_1_io_enq_bits_user;
  wire  Queue_22_1_io_deq_ready;
  wire  Queue_22_1_io_deq_valid;
  wire [1:0] Queue_22_1_io_deq_bits_resp;
  wire [4:0] Queue_22_1_io_deq_bits_id;
  wire  Queue_22_1_io_deq_bits_user;
  wire  Queue_22_1_io_count;
  reg  GEN_1;
  reg [31:0] GEN_3;
  OuterMemorySystem outmemsys (
    .clk(outmemsys_clk),
    .reset(outmemsys_reset),
    .io_tiles_cached_0_acquire_ready(outmemsys_io_tiles_cached_0_acquire_ready),
    .io_tiles_cached_0_acquire_valid(outmemsys_io_tiles_cached_0_acquire_valid),
    .io_tiles_cached_0_acquire_bits_addr_block(outmemsys_io_tiles_cached_0_acquire_bits_addr_block),
    .io_tiles_cached_0_acquire_bits_client_xact_id(outmemsys_io_tiles_cached_0_acquire_bits_client_xact_id),
    .io_tiles_cached_0_acquire_bits_addr_beat(outmemsys_io_tiles_cached_0_acquire_bits_addr_beat),
    .io_tiles_cached_0_acquire_bits_is_builtin_type(outmemsys_io_tiles_cached_0_acquire_bits_is_builtin_type),
    .io_tiles_cached_0_acquire_bits_a_type(outmemsys_io_tiles_cached_0_acquire_bits_a_type),
    .io_tiles_cached_0_acquire_bits_union(outmemsys_io_tiles_cached_0_acquire_bits_union),
    .io_tiles_cached_0_acquire_bits_data(outmemsys_io_tiles_cached_0_acquire_bits_data),
    .io_tiles_cached_0_probe_ready(outmemsys_io_tiles_cached_0_probe_ready),
    .io_tiles_cached_0_probe_valid(outmemsys_io_tiles_cached_0_probe_valid),
    .io_tiles_cached_0_probe_bits_addr_block(outmemsys_io_tiles_cached_0_probe_bits_addr_block),
    .io_tiles_cached_0_probe_bits_p_type(outmemsys_io_tiles_cached_0_probe_bits_p_type),
    .io_tiles_cached_0_release_ready(outmemsys_io_tiles_cached_0_release_ready),
    .io_tiles_cached_0_release_valid(outmemsys_io_tiles_cached_0_release_valid),
    .io_tiles_cached_0_release_bits_addr_beat(outmemsys_io_tiles_cached_0_release_bits_addr_beat),
    .io_tiles_cached_0_release_bits_addr_block(outmemsys_io_tiles_cached_0_release_bits_addr_block),
    .io_tiles_cached_0_release_bits_client_xact_id(outmemsys_io_tiles_cached_0_release_bits_client_xact_id),
    .io_tiles_cached_0_release_bits_voluntary(outmemsys_io_tiles_cached_0_release_bits_voluntary),
    .io_tiles_cached_0_release_bits_r_type(outmemsys_io_tiles_cached_0_release_bits_r_type),
    .io_tiles_cached_0_release_bits_data(outmemsys_io_tiles_cached_0_release_bits_data),
    .io_tiles_cached_0_grant_ready(outmemsys_io_tiles_cached_0_grant_ready),
    .io_tiles_cached_0_grant_valid(outmemsys_io_tiles_cached_0_grant_valid),
    .io_tiles_cached_0_grant_bits_addr_beat(outmemsys_io_tiles_cached_0_grant_bits_addr_beat),
    .io_tiles_cached_0_grant_bits_client_xact_id(outmemsys_io_tiles_cached_0_grant_bits_client_xact_id),
    .io_tiles_cached_0_grant_bits_manager_xact_id(outmemsys_io_tiles_cached_0_grant_bits_manager_xact_id),
    .io_tiles_cached_0_grant_bits_is_builtin_type(outmemsys_io_tiles_cached_0_grant_bits_is_builtin_type),
    .io_tiles_cached_0_grant_bits_g_type(outmemsys_io_tiles_cached_0_grant_bits_g_type),
    .io_tiles_cached_0_grant_bits_data(outmemsys_io_tiles_cached_0_grant_bits_data),
    .io_tiles_cached_0_grant_bits_manager_id(outmemsys_io_tiles_cached_0_grant_bits_manager_id),
    .io_tiles_cached_0_finish_ready(outmemsys_io_tiles_cached_0_finish_ready),
    .io_tiles_cached_0_finish_valid(outmemsys_io_tiles_cached_0_finish_valid),
    .io_tiles_cached_0_finish_bits_manager_xact_id(outmemsys_io_tiles_cached_0_finish_bits_manager_xact_id),
    .io_tiles_cached_0_finish_bits_manager_id(outmemsys_io_tiles_cached_0_finish_bits_manager_id),
    .io_tiles_uncached_0_acquire_ready(outmemsys_io_tiles_uncached_0_acquire_ready),
    .io_tiles_uncached_0_acquire_valid(outmemsys_io_tiles_uncached_0_acquire_valid),
    .io_tiles_uncached_0_acquire_bits_addr_block(outmemsys_io_tiles_uncached_0_acquire_bits_addr_block),
    .io_tiles_uncached_0_acquire_bits_client_xact_id(outmemsys_io_tiles_uncached_0_acquire_bits_client_xact_id),
    .io_tiles_uncached_0_acquire_bits_addr_beat(outmemsys_io_tiles_uncached_0_acquire_bits_addr_beat),
    .io_tiles_uncached_0_acquire_bits_is_builtin_type(outmemsys_io_tiles_uncached_0_acquire_bits_is_builtin_type),
    .io_tiles_uncached_0_acquire_bits_a_type(outmemsys_io_tiles_uncached_0_acquire_bits_a_type),
    .io_tiles_uncached_0_acquire_bits_union(outmemsys_io_tiles_uncached_0_acquire_bits_union),
    .io_tiles_uncached_0_acquire_bits_data(outmemsys_io_tiles_uncached_0_acquire_bits_data),
    .io_tiles_uncached_0_grant_ready(outmemsys_io_tiles_uncached_0_grant_ready),
    .io_tiles_uncached_0_grant_valid(outmemsys_io_tiles_uncached_0_grant_valid),
    .io_tiles_uncached_0_grant_bits_addr_beat(outmemsys_io_tiles_uncached_0_grant_bits_addr_beat),
    .io_tiles_uncached_0_grant_bits_client_xact_id(outmemsys_io_tiles_uncached_0_grant_bits_client_xact_id),
    .io_tiles_uncached_0_grant_bits_manager_xact_id(outmemsys_io_tiles_uncached_0_grant_bits_manager_xact_id),
    .io_tiles_uncached_0_grant_bits_is_builtin_type(outmemsys_io_tiles_uncached_0_grant_bits_is_builtin_type),
    .io_tiles_uncached_0_grant_bits_g_type(outmemsys_io_tiles_uncached_0_grant_bits_g_type),
    .io_tiles_uncached_0_grant_bits_data(outmemsys_io_tiles_uncached_0_grant_bits_data),
    .io_incoherent_0(outmemsys_io_incoherent_0),
    .io_mem_axi_0_aw_ready(outmemsys_io_mem_axi_0_aw_ready),
    .io_mem_axi_0_aw_valid(outmemsys_io_mem_axi_0_aw_valid),
    .io_mem_axi_0_aw_bits_addr(outmemsys_io_mem_axi_0_aw_bits_addr),
    .io_mem_axi_0_aw_bits_len(outmemsys_io_mem_axi_0_aw_bits_len),
    .io_mem_axi_0_aw_bits_size(outmemsys_io_mem_axi_0_aw_bits_size),
    .io_mem_axi_0_aw_bits_burst(outmemsys_io_mem_axi_0_aw_bits_burst),
    .io_mem_axi_0_aw_bits_lock(outmemsys_io_mem_axi_0_aw_bits_lock),
    .io_mem_axi_0_aw_bits_cache(outmemsys_io_mem_axi_0_aw_bits_cache),
    .io_mem_axi_0_aw_bits_prot(outmemsys_io_mem_axi_0_aw_bits_prot),
    .io_mem_axi_0_aw_bits_qos(outmemsys_io_mem_axi_0_aw_bits_qos),
    .io_mem_axi_0_aw_bits_region(outmemsys_io_mem_axi_0_aw_bits_region),
    .io_mem_axi_0_aw_bits_id(outmemsys_io_mem_axi_0_aw_bits_id),
    .io_mem_axi_0_aw_bits_user(outmemsys_io_mem_axi_0_aw_bits_user),
    .io_mem_axi_0_w_ready(outmemsys_io_mem_axi_0_w_ready),
    .io_mem_axi_0_w_valid(outmemsys_io_mem_axi_0_w_valid),
    .io_mem_axi_0_w_bits_data(outmemsys_io_mem_axi_0_w_bits_data),
    .io_mem_axi_0_w_bits_last(outmemsys_io_mem_axi_0_w_bits_last),
    .io_mem_axi_0_w_bits_id(outmemsys_io_mem_axi_0_w_bits_id),
    .io_mem_axi_0_w_bits_strb(outmemsys_io_mem_axi_0_w_bits_strb),
    .io_mem_axi_0_w_bits_user(outmemsys_io_mem_axi_0_w_bits_user),
    .io_mem_axi_0_b_ready(outmemsys_io_mem_axi_0_b_ready),
    .io_mem_axi_0_b_valid(outmemsys_io_mem_axi_0_b_valid),
    .io_mem_axi_0_b_bits_resp(outmemsys_io_mem_axi_0_b_bits_resp),
    .io_mem_axi_0_b_bits_id(outmemsys_io_mem_axi_0_b_bits_id),
    .io_mem_axi_0_b_bits_user(outmemsys_io_mem_axi_0_b_bits_user),
    .io_mem_axi_0_ar_ready(outmemsys_io_mem_axi_0_ar_ready),
    .io_mem_axi_0_ar_valid(outmemsys_io_mem_axi_0_ar_valid),
    .io_mem_axi_0_ar_bits_addr(outmemsys_io_mem_axi_0_ar_bits_addr),
    .io_mem_axi_0_ar_bits_len(outmemsys_io_mem_axi_0_ar_bits_len),
    .io_mem_axi_0_ar_bits_size(outmemsys_io_mem_axi_0_ar_bits_size),
    .io_mem_axi_0_ar_bits_burst(outmemsys_io_mem_axi_0_ar_bits_burst),
    .io_mem_axi_0_ar_bits_lock(outmemsys_io_mem_axi_0_ar_bits_lock),
    .io_mem_axi_0_ar_bits_cache(outmemsys_io_mem_axi_0_ar_bits_cache),
    .io_mem_axi_0_ar_bits_prot(outmemsys_io_mem_axi_0_ar_bits_prot),
    .io_mem_axi_0_ar_bits_qos(outmemsys_io_mem_axi_0_ar_bits_qos),
    .io_mem_axi_0_ar_bits_region(outmemsys_io_mem_axi_0_ar_bits_region),
    .io_mem_axi_0_ar_bits_id(outmemsys_io_mem_axi_0_ar_bits_id),
    .io_mem_axi_0_ar_bits_user(outmemsys_io_mem_axi_0_ar_bits_user),
    .io_mem_axi_0_r_ready(outmemsys_io_mem_axi_0_r_ready),
    .io_mem_axi_0_r_valid(outmemsys_io_mem_axi_0_r_valid),
    .io_mem_axi_0_r_bits_resp(outmemsys_io_mem_axi_0_r_bits_resp),
    .io_mem_axi_0_r_bits_data(outmemsys_io_mem_axi_0_r_bits_data),
    .io_mem_axi_0_r_bits_last(outmemsys_io_mem_axi_0_r_bits_last),
    .io_mem_axi_0_r_bits_id(outmemsys_io_mem_axi_0_r_bits_id),
    .io_mem_axi_0_r_bits_user(outmemsys_io_mem_axi_0_r_bits_user),
    .io_mmio_acquire_ready(outmemsys_io_mmio_acquire_ready),
    .io_mmio_acquire_valid(outmemsys_io_mmio_acquire_valid),
    .io_mmio_acquire_bits_addr_block(outmemsys_io_mmio_acquire_bits_addr_block),
    .io_mmio_acquire_bits_client_xact_id(outmemsys_io_mmio_acquire_bits_client_xact_id),
    .io_mmio_acquire_bits_addr_beat(outmemsys_io_mmio_acquire_bits_addr_beat),
    .io_mmio_acquire_bits_is_builtin_type(outmemsys_io_mmio_acquire_bits_is_builtin_type),
    .io_mmio_acquire_bits_a_type(outmemsys_io_mmio_acquire_bits_a_type),
    .io_mmio_acquire_bits_union(outmemsys_io_mmio_acquire_bits_union),
    .io_mmio_acquire_bits_data(outmemsys_io_mmio_acquire_bits_data),
    .io_mmio_grant_ready(outmemsys_io_mmio_grant_ready),
    .io_mmio_grant_valid(outmemsys_io_mmio_grant_valid),
    .io_mmio_grant_bits_addr_beat(outmemsys_io_mmio_grant_bits_addr_beat),
    .io_mmio_grant_bits_client_xact_id(outmemsys_io_mmio_grant_bits_client_xact_id),
    .io_mmio_grant_bits_manager_xact_id(outmemsys_io_mmio_grant_bits_manager_xact_id),
    .io_mmio_grant_bits_is_builtin_type(outmemsys_io_mmio_grant_bits_is_builtin_type),
    .io_mmio_grant_bits_g_type(outmemsys_io_mmio_grant_bits_g_type),
    .io_mmio_grant_bits_data(outmemsys_io_mmio_grant_bits_data)
  );
  TileLinkRecursiveInterconnect TileLinkRecursiveInterconnect_2 (
    .clk(TileLinkRecursiveInterconnect_2_clk),
    .reset(TileLinkRecursiveInterconnect_2_reset),
    .io_in_0_acquire_ready(TileLinkRecursiveInterconnect_2_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(TileLinkRecursiveInterconnect_2_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(TileLinkRecursiveInterconnect_2_io_in_0_grant_ready),
    .io_in_0_grant_valid(TileLinkRecursiveInterconnect_2_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(TileLinkRecursiveInterconnect_2_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(TileLinkRecursiveInterconnect_2_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(TileLinkRecursiveInterconnect_2_io_out_0_grant_ready),
    .io_out_0_grant_valid(TileLinkRecursiveInterconnect_2_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(TileLinkRecursiveInterconnect_2_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(TileLinkRecursiveInterconnect_2_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(TileLinkRecursiveInterconnect_2_io_out_1_grant_ready),
    .io_out_1_grant_valid(TileLinkRecursiveInterconnect_2_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_data),
    .io_out_2_acquire_ready(TileLinkRecursiveInterconnect_2_io_out_2_acquire_ready),
    .io_out_2_acquire_valid(TileLinkRecursiveInterconnect_2_io_out_2_acquire_valid),
    .io_out_2_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_block),
    .io_out_2_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_client_xact_id),
    .io_out_2_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_beat),
    .io_out_2_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_is_builtin_type),
    .io_out_2_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_a_type),
    .io_out_2_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_union),
    .io_out_2_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_data),
    .io_out_2_grant_ready(TileLinkRecursiveInterconnect_2_io_out_2_grant_ready),
    .io_out_2_grant_valid(TileLinkRecursiveInterconnect_2_io_out_2_grant_valid),
    .io_out_2_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_addr_beat),
    .io_out_2_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_client_xact_id),
    .io_out_2_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_manager_xact_id),
    .io_out_2_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_is_builtin_type),
    .io_out_2_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_g_type),
    .io_out_2_grant_bits_data(TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_data),
    .io_out_3_acquire_ready(TileLinkRecursiveInterconnect_2_io_out_3_acquire_ready),
    .io_out_3_acquire_valid(TileLinkRecursiveInterconnect_2_io_out_3_acquire_valid),
    .io_out_3_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_block),
    .io_out_3_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_client_xact_id),
    .io_out_3_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_beat),
    .io_out_3_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_is_builtin_type),
    .io_out_3_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_a_type),
    .io_out_3_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_union),
    .io_out_3_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_data),
    .io_out_3_grant_ready(TileLinkRecursiveInterconnect_2_io_out_3_grant_ready),
    .io_out_3_grant_valid(TileLinkRecursiveInterconnect_2_io_out_3_grant_valid),
    .io_out_3_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_addr_beat),
    .io_out_3_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_client_xact_id),
    .io_out_3_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_manager_xact_id),
    .io_out_3_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_is_builtin_type),
    .io_out_3_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_g_type),
    .io_out_3_grant_bits_data(TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_data),
    .io_out_4_acquire_ready(TileLinkRecursiveInterconnect_2_io_out_4_acquire_ready),
    .io_out_4_acquire_valid(TileLinkRecursiveInterconnect_2_io_out_4_acquire_valid),
    .io_out_4_acquire_bits_addr_block(TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_addr_block),
    .io_out_4_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_client_xact_id),
    .io_out_4_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_addr_beat),
    .io_out_4_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_is_builtin_type),
    .io_out_4_acquire_bits_a_type(TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_a_type),
    .io_out_4_acquire_bits_union(TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_union),
    .io_out_4_acquire_bits_data(TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_data),
    .io_out_4_grant_ready(TileLinkRecursiveInterconnect_2_io_out_4_grant_ready),
    .io_out_4_grant_valid(TileLinkRecursiveInterconnect_2_io_out_4_grant_valid),
    .io_out_4_grant_bits_addr_beat(TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_addr_beat),
    .io_out_4_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_client_xact_id),
    .io_out_4_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_manager_xact_id),
    .io_out_4_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_is_builtin_type),
    .io_out_4_grant_bits_g_type(TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_g_type),
    .io_out_4_grant_bits_data(TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_data)
  );
  PLIC PLIC_1 (
    .clk(PLIC_1_clk),
    .reset(PLIC_1_reset),
    .io_devices_0_valid(PLIC_1_io_devices_0_valid),
    .io_devices_0_ready(PLIC_1_io_devices_0_ready),
    .io_devices_0_complete(PLIC_1_io_devices_0_complete),
    .io_devices_1_valid(PLIC_1_io_devices_1_valid),
    .io_devices_1_ready(PLIC_1_io_devices_1_ready),
    .io_devices_1_complete(PLIC_1_io_devices_1_complete),
    .io_devices_2_valid(PLIC_1_io_devices_2_valid),
    .io_devices_2_ready(PLIC_1_io_devices_2_ready),
    .io_devices_2_complete(PLIC_1_io_devices_2_complete),
    .io_devices_3_valid(PLIC_1_io_devices_3_valid),
    .io_devices_3_ready(PLIC_1_io_devices_3_ready),
    .io_devices_3_complete(PLIC_1_io_devices_3_complete),
    .io_devices_4_valid(PLIC_1_io_devices_4_valid),
    .io_devices_4_ready(PLIC_1_io_devices_4_ready),
    .io_devices_4_complete(PLIC_1_io_devices_4_complete),
    .io_devices_5_valid(PLIC_1_io_devices_5_valid),
    .io_devices_5_ready(PLIC_1_io_devices_5_ready),
    .io_devices_5_complete(PLIC_1_io_devices_5_complete),
    .io_devices_6_valid(PLIC_1_io_devices_6_valid),
    .io_devices_6_ready(PLIC_1_io_devices_6_ready),
    .io_devices_6_complete(PLIC_1_io_devices_6_complete),
    .io_devices_7_valid(PLIC_1_io_devices_7_valid),
    .io_devices_7_ready(PLIC_1_io_devices_7_ready),
    .io_devices_7_complete(PLIC_1_io_devices_7_complete),
    .io_devices_8_valid(PLIC_1_io_devices_8_valid),
    .io_devices_8_ready(PLIC_1_io_devices_8_ready),
    .io_devices_8_complete(PLIC_1_io_devices_8_complete),
    .io_devices_9_valid(PLIC_1_io_devices_9_valid),
    .io_devices_9_ready(PLIC_1_io_devices_9_ready),
    .io_devices_9_complete(PLIC_1_io_devices_9_complete),
    .io_devices_10_valid(PLIC_1_io_devices_10_valid),
    .io_devices_10_ready(PLIC_1_io_devices_10_ready),
    .io_devices_10_complete(PLIC_1_io_devices_10_complete),
    .io_devices_11_valid(PLIC_1_io_devices_11_valid),
    .io_devices_11_ready(PLIC_1_io_devices_11_ready),
    .io_devices_11_complete(PLIC_1_io_devices_11_complete),
    .io_devices_12_valid(PLIC_1_io_devices_12_valid),
    .io_devices_12_ready(PLIC_1_io_devices_12_ready),
    .io_devices_12_complete(PLIC_1_io_devices_12_complete),
    .io_devices_13_valid(PLIC_1_io_devices_13_valid),
    .io_devices_13_ready(PLIC_1_io_devices_13_ready),
    .io_devices_13_complete(PLIC_1_io_devices_13_complete),
    .io_devices_14_valid(PLIC_1_io_devices_14_valid),
    .io_devices_14_ready(PLIC_1_io_devices_14_ready),
    .io_devices_14_complete(PLIC_1_io_devices_14_complete),
    .io_devices_15_valid(PLIC_1_io_devices_15_valid),
    .io_devices_15_ready(PLIC_1_io_devices_15_ready),
    .io_devices_15_complete(PLIC_1_io_devices_15_complete),
    .io_devices_16_valid(PLIC_1_io_devices_16_valid),
    .io_devices_16_ready(PLIC_1_io_devices_16_ready),
    .io_devices_16_complete(PLIC_1_io_devices_16_complete),
    .io_devices_17_valid(PLIC_1_io_devices_17_valid),
    .io_devices_17_ready(PLIC_1_io_devices_17_ready),
    .io_devices_17_complete(PLIC_1_io_devices_17_complete),
    .io_devices_18_valid(PLIC_1_io_devices_18_valid),
    .io_devices_18_ready(PLIC_1_io_devices_18_ready),
    .io_devices_18_complete(PLIC_1_io_devices_18_complete),
    .io_devices_19_valid(PLIC_1_io_devices_19_valid),
    .io_devices_19_ready(PLIC_1_io_devices_19_ready),
    .io_devices_19_complete(PLIC_1_io_devices_19_complete),
    .io_devices_20_valid(PLIC_1_io_devices_20_valid),
    .io_devices_20_ready(PLIC_1_io_devices_20_ready),
    .io_devices_20_complete(PLIC_1_io_devices_20_complete),
    .io_devices_21_valid(PLIC_1_io_devices_21_valid),
    .io_devices_21_ready(PLIC_1_io_devices_21_ready),
    .io_devices_21_complete(PLIC_1_io_devices_21_complete),
    .io_devices_22_valid(PLIC_1_io_devices_22_valid),
    .io_devices_22_ready(PLIC_1_io_devices_22_ready),
    .io_devices_22_complete(PLIC_1_io_devices_22_complete),
    .io_devices_23_valid(PLIC_1_io_devices_23_valid),
    .io_devices_23_ready(PLIC_1_io_devices_23_ready),
    .io_devices_23_complete(PLIC_1_io_devices_23_complete),
    .io_devices_24_valid(PLIC_1_io_devices_24_valid),
    .io_devices_24_ready(PLIC_1_io_devices_24_ready),
    .io_devices_24_complete(PLIC_1_io_devices_24_complete),
    .io_devices_25_valid(PLIC_1_io_devices_25_valid),
    .io_devices_25_ready(PLIC_1_io_devices_25_ready),
    .io_devices_25_complete(PLIC_1_io_devices_25_complete),
    .io_devices_26_valid(PLIC_1_io_devices_26_valid),
    .io_devices_26_ready(PLIC_1_io_devices_26_ready),
    .io_devices_26_complete(PLIC_1_io_devices_26_complete),
    .io_devices_27_valid(PLIC_1_io_devices_27_valid),
    .io_devices_27_ready(PLIC_1_io_devices_27_ready),
    .io_devices_27_complete(PLIC_1_io_devices_27_complete),
    .io_devices_28_valid(PLIC_1_io_devices_28_valid),
    .io_devices_28_ready(PLIC_1_io_devices_28_ready),
    .io_devices_28_complete(PLIC_1_io_devices_28_complete),
    .io_devices_29_valid(PLIC_1_io_devices_29_valid),
    .io_devices_29_ready(PLIC_1_io_devices_29_ready),
    .io_devices_29_complete(PLIC_1_io_devices_29_complete),
    .io_devices_30_valid(PLIC_1_io_devices_30_valid),
    .io_devices_30_ready(PLIC_1_io_devices_30_ready),
    .io_devices_30_complete(PLIC_1_io_devices_30_complete),
    .io_harts_0(PLIC_1_io_harts_0),
    .io_tl_acquire_ready(PLIC_1_io_tl_acquire_ready),
    .io_tl_acquire_valid(PLIC_1_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(PLIC_1_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(PLIC_1_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(PLIC_1_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(PLIC_1_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(PLIC_1_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(PLIC_1_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(PLIC_1_io_tl_acquire_bits_data),
    .io_tl_grant_ready(PLIC_1_io_tl_grant_ready),
    .io_tl_grant_valid(PLIC_1_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(PLIC_1_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(PLIC_1_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(PLIC_1_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(PLIC_1_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(PLIC_1_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(PLIC_1_io_tl_grant_bits_data)
  );
  LevelGateway LevelGateway_31 (
    .clk(LevelGateway_31_clk),
    .reset(LevelGateway_31_reset),
    .io_interrupt(LevelGateway_31_io_interrupt),
    .io_plic_valid(LevelGateway_31_io_plic_valid),
    .io_plic_ready(LevelGateway_31_io_plic_ready),
    .io_plic_complete(LevelGateway_31_io_plic_complete)
  );
  LevelGateway LevelGateway_1_1 (
    .clk(LevelGateway_1_1_clk),
    .reset(LevelGateway_1_1_reset),
    .io_interrupt(LevelGateway_1_1_io_interrupt),
    .io_plic_valid(LevelGateway_1_1_io_plic_valid),
    .io_plic_ready(LevelGateway_1_1_io_plic_ready),
    .io_plic_complete(LevelGateway_1_1_io_plic_complete)
  );
  LevelGateway LevelGateway_2_1 (
    .clk(LevelGateway_2_1_clk),
    .reset(LevelGateway_2_1_reset),
    .io_interrupt(LevelGateway_2_1_io_interrupt),
    .io_plic_valid(LevelGateway_2_1_io_plic_valid),
    .io_plic_ready(LevelGateway_2_1_io_plic_ready),
    .io_plic_complete(LevelGateway_2_1_io_plic_complete)
  );
  LevelGateway LevelGateway_3_1 (
    .clk(LevelGateway_3_1_clk),
    .reset(LevelGateway_3_1_reset),
    .io_interrupt(LevelGateway_3_1_io_interrupt),
    .io_plic_valid(LevelGateway_3_1_io_plic_valid),
    .io_plic_ready(LevelGateway_3_1_io_plic_ready),
    .io_plic_complete(LevelGateway_3_1_io_plic_complete)
  );
  LevelGateway LevelGateway_4_1 (
    .clk(LevelGateway_4_1_clk),
    .reset(LevelGateway_4_1_reset),
    .io_interrupt(LevelGateway_4_1_io_interrupt),
    .io_plic_valid(LevelGateway_4_1_io_plic_valid),
    .io_plic_ready(LevelGateway_4_1_io_plic_ready),
    .io_plic_complete(LevelGateway_4_1_io_plic_complete)
  );
  LevelGateway LevelGateway_5_1 (
    .clk(LevelGateway_5_1_clk),
    .reset(LevelGateway_5_1_reset),
    .io_interrupt(LevelGateway_5_1_io_interrupt),
    .io_plic_valid(LevelGateway_5_1_io_plic_valid),
    .io_plic_ready(LevelGateway_5_1_io_plic_ready),
    .io_plic_complete(LevelGateway_5_1_io_plic_complete)
  );
  LevelGateway LevelGateway_6_1 (
    .clk(LevelGateway_6_1_clk),
    .reset(LevelGateway_6_1_reset),
    .io_interrupt(LevelGateway_6_1_io_interrupt),
    .io_plic_valid(LevelGateway_6_1_io_plic_valid),
    .io_plic_ready(LevelGateway_6_1_io_plic_ready),
    .io_plic_complete(LevelGateway_6_1_io_plic_complete)
  );
  LevelGateway LevelGateway_7_1 (
    .clk(LevelGateway_7_1_clk),
    .reset(LevelGateway_7_1_reset),
    .io_interrupt(LevelGateway_7_1_io_interrupt),
    .io_plic_valid(LevelGateway_7_1_io_plic_valid),
    .io_plic_ready(LevelGateway_7_1_io_plic_ready),
    .io_plic_complete(LevelGateway_7_1_io_plic_complete)
  );
  LevelGateway LevelGateway_8_1 (
    .clk(LevelGateway_8_1_clk),
    .reset(LevelGateway_8_1_reset),
    .io_interrupt(LevelGateway_8_1_io_interrupt),
    .io_plic_valid(LevelGateway_8_1_io_plic_valid),
    .io_plic_ready(LevelGateway_8_1_io_plic_ready),
    .io_plic_complete(LevelGateway_8_1_io_plic_complete)
  );
  LevelGateway LevelGateway_9_1 (
    .clk(LevelGateway_9_1_clk),
    .reset(LevelGateway_9_1_reset),
    .io_interrupt(LevelGateway_9_1_io_interrupt),
    .io_plic_valid(LevelGateway_9_1_io_plic_valid),
    .io_plic_ready(LevelGateway_9_1_io_plic_ready),
    .io_plic_complete(LevelGateway_9_1_io_plic_complete)
  );
  LevelGateway LevelGateway_10_1 (
    .clk(LevelGateway_10_1_clk),
    .reset(LevelGateway_10_1_reset),
    .io_interrupt(LevelGateway_10_1_io_interrupt),
    .io_plic_valid(LevelGateway_10_1_io_plic_valid),
    .io_plic_ready(LevelGateway_10_1_io_plic_ready),
    .io_plic_complete(LevelGateway_10_1_io_plic_complete)
  );
  LevelGateway LevelGateway_11_1 (
    .clk(LevelGateway_11_1_clk),
    .reset(LevelGateway_11_1_reset),
    .io_interrupt(LevelGateway_11_1_io_interrupt),
    .io_plic_valid(LevelGateway_11_1_io_plic_valid),
    .io_plic_ready(LevelGateway_11_1_io_plic_ready),
    .io_plic_complete(LevelGateway_11_1_io_plic_complete)
  );
  LevelGateway LevelGateway_12_1 (
    .clk(LevelGateway_12_1_clk),
    .reset(LevelGateway_12_1_reset),
    .io_interrupt(LevelGateway_12_1_io_interrupt),
    .io_plic_valid(LevelGateway_12_1_io_plic_valid),
    .io_plic_ready(LevelGateway_12_1_io_plic_ready),
    .io_plic_complete(LevelGateway_12_1_io_plic_complete)
  );
  LevelGateway LevelGateway_13_1 (
    .clk(LevelGateway_13_1_clk),
    .reset(LevelGateway_13_1_reset),
    .io_interrupt(LevelGateway_13_1_io_interrupt),
    .io_plic_valid(LevelGateway_13_1_io_plic_valid),
    .io_plic_ready(LevelGateway_13_1_io_plic_ready),
    .io_plic_complete(LevelGateway_13_1_io_plic_complete)
  );
  LevelGateway LevelGateway_14_1 (
    .clk(LevelGateway_14_1_clk),
    .reset(LevelGateway_14_1_reset),
    .io_interrupt(LevelGateway_14_1_io_interrupt),
    .io_plic_valid(LevelGateway_14_1_io_plic_valid),
    .io_plic_ready(LevelGateway_14_1_io_plic_ready),
    .io_plic_complete(LevelGateway_14_1_io_plic_complete)
  );
  LevelGateway LevelGateway_15_1 (
    .clk(LevelGateway_15_1_clk),
    .reset(LevelGateway_15_1_reset),
    .io_interrupt(LevelGateway_15_1_io_interrupt),
    .io_plic_valid(LevelGateway_15_1_io_plic_valid),
    .io_plic_ready(LevelGateway_15_1_io_plic_ready),
    .io_plic_complete(LevelGateway_15_1_io_plic_complete)
  );
  LevelGateway LevelGateway_16_1 (
    .clk(LevelGateway_16_1_clk),
    .reset(LevelGateway_16_1_reset),
    .io_interrupt(LevelGateway_16_1_io_interrupt),
    .io_plic_valid(LevelGateway_16_1_io_plic_valid),
    .io_plic_ready(LevelGateway_16_1_io_plic_ready),
    .io_plic_complete(LevelGateway_16_1_io_plic_complete)
  );
  LevelGateway LevelGateway_17_1 (
    .clk(LevelGateway_17_1_clk),
    .reset(LevelGateway_17_1_reset),
    .io_interrupt(LevelGateway_17_1_io_interrupt),
    .io_plic_valid(LevelGateway_17_1_io_plic_valid),
    .io_plic_ready(LevelGateway_17_1_io_plic_ready),
    .io_plic_complete(LevelGateway_17_1_io_plic_complete)
  );
  LevelGateway LevelGateway_18_1 (
    .clk(LevelGateway_18_1_clk),
    .reset(LevelGateway_18_1_reset),
    .io_interrupt(LevelGateway_18_1_io_interrupt),
    .io_plic_valid(LevelGateway_18_1_io_plic_valid),
    .io_plic_ready(LevelGateway_18_1_io_plic_ready),
    .io_plic_complete(LevelGateway_18_1_io_plic_complete)
  );
  LevelGateway LevelGateway_19_1 (
    .clk(LevelGateway_19_1_clk),
    .reset(LevelGateway_19_1_reset),
    .io_interrupt(LevelGateway_19_1_io_interrupt),
    .io_plic_valid(LevelGateway_19_1_io_plic_valid),
    .io_plic_ready(LevelGateway_19_1_io_plic_ready),
    .io_plic_complete(LevelGateway_19_1_io_plic_complete)
  );
  LevelGateway LevelGateway_20_1 (
    .clk(LevelGateway_20_1_clk),
    .reset(LevelGateway_20_1_reset),
    .io_interrupt(LevelGateway_20_1_io_interrupt),
    .io_plic_valid(LevelGateway_20_1_io_plic_valid),
    .io_plic_ready(LevelGateway_20_1_io_plic_ready),
    .io_plic_complete(LevelGateway_20_1_io_plic_complete)
  );
  LevelGateway LevelGateway_21_1 (
    .clk(LevelGateway_21_1_clk),
    .reset(LevelGateway_21_1_reset),
    .io_interrupt(LevelGateway_21_1_io_interrupt),
    .io_plic_valid(LevelGateway_21_1_io_plic_valid),
    .io_plic_ready(LevelGateway_21_1_io_plic_ready),
    .io_plic_complete(LevelGateway_21_1_io_plic_complete)
  );
  LevelGateway LevelGateway_22_1 (
    .clk(LevelGateway_22_1_clk),
    .reset(LevelGateway_22_1_reset),
    .io_interrupt(LevelGateway_22_1_io_interrupt),
    .io_plic_valid(LevelGateway_22_1_io_plic_valid),
    .io_plic_ready(LevelGateway_22_1_io_plic_ready),
    .io_plic_complete(LevelGateway_22_1_io_plic_complete)
  );
  LevelGateway LevelGateway_23_1 (
    .clk(LevelGateway_23_1_clk),
    .reset(LevelGateway_23_1_reset),
    .io_interrupt(LevelGateway_23_1_io_interrupt),
    .io_plic_valid(LevelGateway_23_1_io_plic_valid),
    .io_plic_ready(LevelGateway_23_1_io_plic_ready),
    .io_plic_complete(LevelGateway_23_1_io_plic_complete)
  );
  LevelGateway LevelGateway_24_1 (
    .clk(LevelGateway_24_1_clk),
    .reset(LevelGateway_24_1_reset),
    .io_interrupt(LevelGateway_24_1_io_interrupt),
    .io_plic_valid(LevelGateway_24_1_io_plic_valid),
    .io_plic_ready(LevelGateway_24_1_io_plic_ready),
    .io_plic_complete(LevelGateway_24_1_io_plic_complete)
  );
  LevelGateway LevelGateway_25_1 (
    .clk(LevelGateway_25_1_clk),
    .reset(LevelGateway_25_1_reset),
    .io_interrupt(LevelGateway_25_1_io_interrupt),
    .io_plic_valid(LevelGateway_25_1_io_plic_valid),
    .io_plic_ready(LevelGateway_25_1_io_plic_ready),
    .io_plic_complete(LevelGateway_25_1_io_plic_complete)
  );
  LevelGateway LevelGateway_26_1 (
    .clk(LevelGateway_26_1_clk),
    .reset(LevelGateway_26_1_reset),
    .io_interrupt(LevelGateway_26_1_io_interrupt),
    .io_plic_valid(LevelGateway_26_1_io_plic_valid),
    .io_plic_ready(LevelGateway_26_1_io_plic_ready),
    .io_plic_complete(LevelGateway_26_1_io_plic_complete)
  );
  LevelGateway LevelGateway_27_1 (
    .clk(LevelGateway_27_1_clk),
    .reset(LevelGateway_27_1_reset),
    .io_interrupt(LevelGateway_27_1_io_interrupt),
    .io_plic_valid(LevelGateway_27_1_io_plic_valid),
    .io_plic_ready(LevelGateway_27_1_io_plic_ready),
    .io_plic_complete(LevelGateway_27_1_io_plic_complete)
  );
  LevelGateway LevelGateway_28_1 (
    .clk(LevelGateway_28_1_clk),
    .reset(LevelGateway_28_1_reset),
    .io_interrupt(LevelGateway_28_1_io_interrupt),
    .io_plic_valid(LevelGateway_28_1_io_plic_valid),
    .io_plic_ready(LevelGateway_28_1_io_plic_ready),
    .io_plic_complete(LevelGateway_28_1_io_plic_complete)
  );
  LevelGateway LevelGateway_29_1 (
    .clk(LevelGateway_29_1_clk),
    .reset(LevelGateway_29_1_reset),
    .io_interrupt(LevelGateway_29_1_io_interrupt),
    .io_plic_valid(LevelGateway_29_1_io_plic_valid),
    .io_plic_ready(LevelGateway_29_1_io_plic_ready),
    .io_plic_complete(LevelGateway_29_1_io_plic_complete)
  );
  LevelGateway LevelGateway_30_1 (
    .clk(LevelGateway_30_1_clk),
    .reset(LevelGateway_30_1_reset),
    .io_interrupt(LevelGateway_30_1_io_interrupt),
    .io_plic_valid(LevelGateway_30_1_io_plic_valid),
    .io_plic_ready(LevelGateway_30_1_io_plic_ready),
    .io_plic_complete(LevelGateway_30_1_io_plic_complete)
  );
  DebugModule DebugModule_1 (
    .clk(DebugModule_1_clk),
    .reset(DebugModule_1_reset),
    .io_db_req_ready(DebugModule_1_io_db_req_ready),
    .io_db_req_valid(DebugModule_1_io_db_req_valid),
    .io_db_req_bits_addr(DebugModule_1_io_db_req_bits_addr),
    .io_db_req_bits_op(DebugModule_1_io_db_req_bits_op),
    .io_db_req_bits_data(DebugModule_1_io_db_req_bits_data),
    .io_db_resp_ready(DebugModule_1_io_db_resp_ready),
    .io_db_resp_valid(DebugModule_1_io_db_resp_valid),
    .io_db_resp_bits_resp(DebugModule_1_io_db_resp_bits_resp),
    .io_db_resp_bits_data(DebugModule_1_io_db_resp_bits_data),
    .io_debugInterrupts_0(DebugModule_1_io_debugInterrupts_0),
    .io_tl_acquire_ready(DebugModule_1_io_tl_acquire_ready),
    .io_tl_acquire_valid(DebugModule_1_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(DebugModule_1_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(DebugModule_1_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(DebugModule_1_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(DebugModule_1_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(DebugModule_1_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(DebugModule_1_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(DebugModule_1_io_tl_acquire_bits_data),
    .io_tl_grant_ready(DebugModule_1_io_tl_grant_ready),
    .io_tl_grant_valid(DebugModule_1_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(DebugModule_1_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(DebugModule_1_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(DebugModule_1_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(DebugModule_1_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(DebugModule_1_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(DebugModule_1_io_tl_grant_bits_data),
    .io_ndreset(DebugModule_1_io_ndreset),
    .io_fullreset(DebugModule_1_io_fullreset)
  );
  PRCI PRCI_1 (
    .clk(PRCI_1_clk),
    .reset(PRCI_1_reset),
    .io_interrupts_0_meip(PRCI_1_io_interrupts_0_meip),
    .io_interrupts_0_seip(PRCI_1_io_interrupts_0_seip),
    .io_interrupts_0_debug(PRCI_1_io_interrupts_0_debug),
    .io_tl_acquire_ready(PRCI_1_io_tl_acquire_ready),
    .io_tl_acquire_valid(PRCI_1_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(PRCI_1_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(PRCI_1_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(PRCI_1_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(PRCI_1_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(PRCI_1_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(PRCI_1_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(PRCI_1_io_tl_acquire_bits_data),
    .io_tl_grant_ready(PRCI_1_io_tl_grant_ready),
    .io_tl_grant_valid(PRCI_1_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(PRCI_1_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(PRCI_1_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(PRCI_1_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(PRCI_1_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(PRCI_1_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(PRCI_1_io_tl_grant_bits_data),
    .io_tiles_0_reset(PRCI_1_io_tiles_0_reset),
    .io_tiles_0_id(PRCI_1_io_tiles_0_id),
    .io_tiles_0_interrupts_meip(PRCI_1_io_tiles_0_interrupts_meip),
    .io_tiles_0_interrupts_seip(PRCI_1_io_tiles_0_interrupts_seip),
    .io_tiles_0_interrupts_debug(PRCI_1_io_tiles_0_interrupts_debug),
    .io_tiles_0_interrupts_mtip(PRCI_1_io_tiles_0_interrupts_mtip),
    .io_tiles_0_interrupts_msip(PRCI_1_io_tiles_0_interrupts_msip),
    .io_rtcTick(PRCI_1_io_rtcTick)
  );
  ROMSlave ROMSlave_1 (
    .clk(ROMSlave_1_clk),
    .reset(ROMSlave_1_reset),
    .io_acquire_ready(ROMSlave_1_io_acquire_ready),
    .io_acquire_valid(ROMSlave_1_io_acquire_valid),
    .io_acquire_bits_addr_block(ROMSlave_1_io_acquire_bits_addr_block),
    .io_acquire_bits_client_xact_id(ROMSlave_1_io_acquire_bits_client_xact_id),
    .io_acquire_bits_addr_beat(ROMSlave_1_io_acquire_bits_addr_beat),
    .io_acquire_bits_is_builtin_type(ROMSlave_1_io_acquire_bits_is_builtin_type),
    .io_acquire_bits_a_type(ROMSlave_1_io_acquire_bits_a_type),
    .io_acquire_bits_union(ROMSlave_1_io_acquire_bits_union),
    .io_acquire_bits_data(ROMSlave_1_io_acquire_bits_data),
    .io_grant_ready(ROMSlave_1_io_grant_ready),
    .io_grant_valid(ROMSlave_1_io_grant_valid),
    .io_grant_bits_addr_beat(ROMSlave_1_io_grant_bits_addr_beat),
    .io_grant_bits_client_xact_id(ROMSlave_1_io_grant_bits_client_xact_id),
    .io_grant_bits_manager_xact_id(ROMSlave_1_io_grant_bits_manager_xact_id),
    .io_grant_bits_is_builtin_type(ROMSlave_1_io_grant_bits_is_builtin_type),
    .io_grant_bits_g_type(ROMSlave_1_io_grant_bits_g_type),
    .io_grant_bits_data(ROMSlave_1_io_grant_bits_data)
  );
  NastiIOTileLinkIOConverter_1 NastiIOTileLinkIOConverter_1_1 (
    .clk(NastiIOTileLinkIOConverter_1_1_clk),
    .reset(NastiIOTileLinkIOConverter_1_1_reset),
    .io_tl_acquire_ready(NastiIOTileLinkIOConverter_1_1_io_tl_acquire_ready),
    .io_tl_acquire_valid(NastiIOTileLinkIOConverter_1_1_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_data),
    .io_tl_grant_ready(NastiIOTileLinkIOConverter_1_1_io_tl_grant_ready),
    .io_tl_grant_valid(NastiIOTileLinkIOConverter_1_1_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_data),
    .io_nasti_aw_ready(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_ready),
    .io_nasti_aw_valid(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_valid),
    .io_nasti_aw_bits_addr(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_addr),
    .io_nasti_aw_bits_len(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_len),
    .io_nasti_aw_bits_size(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_size),
    .io_nasti_aw_bits_burst(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_burst),
    .io_nasti_aw_bits_lock(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_lock),
    .io_nasti_aw_bits_cache(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_cache),
    .io_nasti_aw_bits_prot(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_prot),
    .io_nasti_aw_bits_qos(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_qos),
    .io_nasti_aw_bits_region(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_region),
    .io_nasti_aw_bits_id(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_id),
    .io_nasti_aw_bits_user(NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_user),
    .io_nasti_w_ready(NastiIOTileLinkIOConverter_1_1_io_nasti_w_ready),
    .io_nasti_w_valid(NastiIOTileLinkIOConverter_1_1_io_nasti_w_valid),
    .io_nasti_w_bits_data(NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_data),
    .io_nasti_w_bits_last(NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_last),
    .io_nasti_w_bits_id(NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_id),
    .io_nasti_w_bits_strb(NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_strb),
    .io_nasti_w_bits_user(NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_user),
    .io_nasti_b_ready(NastiIOTileLinkIOConverter_1_1_io_nasti_b_ready),
    .io_nasti_b_valid(NastiIOTileLinkIOConverter_1_1_io_nasti_b_valid),
    .io_nasti_b_bits_resp(NastiIOTileLinkIOConverter_1_1_io_nasti_b_bits_resp),
    .io_nasti_b_bits_id(NastiIOTileLinkIOConverter_1_1_io_nasti_b_bits_id),
    .io_nasti_b_bits_user(NastiIOTileLinkIOConverter_1_1_io_nasti_b_bits_user),
    .io_nasti_ar_ready(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_ready),
    .io_nasti_ar_valid(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_valid),
    .io_nasti_ar_bits_addr(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_addr),
    .io_nasti_ar_bits_len(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_len),
    .io_nasti_ar_bits_size(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_size),
    .io_nasti_ar_bits_burst(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_burst),
    .io_nasti_ar_bits_lock(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_lock),
    .io_nasti_ar_bits_cache(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_cache),
    .io_nasti_ar_bits_prot(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_prot),
    .io_nasti_ar_bits_qos(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_qos),
    .io_nasti_ar_bits_region(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_region),
    .io_nasti_ar_bits_id(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_id),
    .io_nasti_ar_bits_user(NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_user),
    .io_nasti_r_ready(NastiIOTileLinkIOConverter_1_1_io_nasti_r_ready),
    .io_nasti_r_valid(NastiIOTileLinkIOConverter_1_1_io_nasti_r_valid),
    .io_nasti_r_bits_resp(NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_resp),
    .io_nasti_r_bits_data(NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_data),
    .io_nasti_r_bits_last(NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_last),
    .io_nasti_r_bits_id(NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_id),
    .io_nasti_r_bits_user(NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_user)
  );
  Queue_10 Queue_18_1 (
    .clk(Queue_18_1_clk),
    .reset(Queue_18_1_reset),
    .io_enq_ready(Queue_18_1_io_enq_ready),
    .io_enq_valid(Queue_18_1_io_enq_valid),
    .io_enq_bits_addr(Queue_18_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_18_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_18_1_io_enq_bits_size),
    .io_enq_bits_burst(Queue_18_1_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_18_1_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_18_1_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_18_1_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_18_1_io_enq_bits_qos),
    .io_enq_bits_region(Queue_18_1_io_enq_bits_region),
    .io_enq_bits_id(Queue_18_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_18_1_io_enq_bits_user),
    .io_deq_ready(Queue_18_1_io_deq_ready),
    .io_deq_valid(Queue_18_1_io_deq_valid),
    .io_deq_bits_addr(Queue_18_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_18_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_18_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_18_1_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_18_1_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_18_1_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_18_1_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_18_1_io_deq_bits_qos),
    .io_deq_bits_region(Queue_18_1_io_deq_bits_region),
    .io_deq_bits_id(Queue_18_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_18_1_io_deq_bits_user),
    .io_count(Queue_18_1_io_count)
  );
  Queue_10 Queue_19_1 (
    .clk(Queue_19_1_clk),
    .reset(Queue_19_1_reset),
    .io_enq_ready(Queue_19_1_io_enq_ready),
    .io_enq_valid(Queue_19_1_io_enq_valid),
    .io_enq_bits_addr(Queue_19_1_io_enq_bits_addr),
    .io_enq_bits_len(Queue_19_1_io_enq_bits_len),
    .io_enq_bits_size(Queue_19_1_io_enq_bits_size),
    .io_enq_bits_burst(Queue_19_1_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_19_1_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_19_1_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_19_1_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_19_1_io_enq_bits_qos),
    .io_enq_bits_region(Queue_19_1_io_enq_bits_region),
    .io_enq_bits_id(Queue_19_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_19_1_io_enq_bits_user),
    .io_deq_ready(Queue_19_1_io_deq_ready),
    .io_deq_valid(Queue_19_1_io_deq_valid),
    .io_deq_bits_addr(Queue_19_1_io_deq_bits_addr),
    .io_deq_bits_len(Queue_19_1_io_deq_bits_len),
    .io_deq_bits_size(Queue_19_1_io_deq_bits_size),
    .io_deq_bits_burst(Queue_19_1_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_19_1_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_19_1_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_19_1_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_19_1_io_deq_bits_qos),
    .io_deq_bits_region(Queue_19_1_io_deq_bits_region),
    .io_deq_bits_id(Queue_19_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_19_1_io_deq_bits_user),
    .io_count(Queue_19_1_io_count)
  );
  Queue_12 Queue_20_1 (
    .clk(Queue_20_1_clk),
    .reset(Queue_20_1_reset),
    .io_enq_ready(Queue_20_1_io_enq_ready),
    .io_enq_valid(Queue_20_1_io_enq_valid),
    .io_enq_bits_data(Queue_20_1_io_enq_bits_data),
    .io_enq_bits_last(Queue_20_1_io_enq_bits_last),
    .io_enq_bits_id(Queue_20_1_io_enq_bits_id),
    .io_enq_bits_strb(Queue_20_1_io_enq_bits_strb),
    .io_enq_bits_user(Queue_20_1_io_enq_bits_user),
    .io_deq_ready(Queue_20_1_io_deq_ready),
    .io_deq_valid(Queue_20_1_io_deq_valid),
    .io_deq_bits_data(Queue_20_1_io_deq_bits_data),
    .io_deq_bits_last(Queue_20_1_io_deq_bits_last),
    .io_deq_bits_id(Queue_20_1_io_deq_bits_id),
    .io_deq_bits_strb(Queue_20_1_io_deq_bits_strb),
    .io_deq_bits_user(Queue_20_1_io_deq_bits_user),
    .io_count(Queue_20_1_io_count)
  );
  Queue_13 Queue_21_1 (
    .clk(Queue_21_1_clk),
    .reset(Queue_21_1_reset),
    .io_enq_ready(Queue_21_1_io_enq_ready),
    .io_enq_valid(Queue_21_1_io_enq_valid),
    .io_enq_bits_resp(Queue_21_1_io_enq_bits_resp),
    .io_enq_bits_data(Queue_21_1_io_enq_bits_data),
    .io_enq_bits_last(Queue_21_1_io_enq_bits_last),
    .io_enq_bits_id(Queue_21_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_21_1_io_enq_bits_user),
    .io_deq_ready(Queue_21_1_io_deq_ready),
    .io_deq_valid(Queue_21_1_io_deq_valid),
    .io_deq_bits_resp(Queue_21_1_io_deq_bits_resp),
    .io_deq_bits_data(Queue_21_1_io_deq_bits_data),
    .io_deq_bits_last(Queue_21_1_io_deq_bits_last),
    .io_deq_bits_id(Queue_21_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_21_1_io_deq_bits_user),
    .io_count(Queue_21_1_io_count)
  );
  Queue_14 Queue_22_1 (
    .clk(Queue_22_1_clk),
    .reset(Queue_22_1_reset),
    .io_enq_ready(Queue_22_1_io_enq_ready),
    .io_enq_valid(Queue_22_1_io_enq_valid),
    .io_enq_bits_resp(Queue_22_1_io_enq_bits_resp),
    .io_enq_bits_id(Queue_22_1_io_enq_bits_id),
    .io_enq_bits_user(Queue_22_1_io_enq_bits_user),
    .io_deq_ready(Queue_22_1_io_deq_ready),
    .io_deq_valid(Queue_22_1_io_deq_valid),
    .io_deq_bits_resp(Queue_22_1_io_deq_bits_resp),
    .io_deq_bits_id(Queue_22_1_io_deq_bits_id),
    .io_deq_bits_user(Queue_22_1_io_deq_bits_user),
    .io_count(Queue_22_1_io_count)
  );
  assign io_mem_axi_0_aw_valid = outmemsys_io_mem_axi_0_aw_valid;
  assign io_mem_axi_0_aw_bits_addr = outmemsys_io_mem_axi_0_aw_bits_addr;
  assign io_mem_axi_0_aw_bits_len = outmemsys_io_mem_axi_0_aw_bits_len;
  assign io_mem_axi_0_aw_bits_size = outmemsys_io_mem_axi_0_aw_bits_size;
  assign io_mem_axi_0_aw_bits_burst = outmemsys_io_mem_axi_0_aw_bits_burst;
  assign io_mem_axi_0_aw_bits_lock = outmemsys_io_mem_axi_0_aw_bits_lock;
  assign io_mem_axi_0_aw_bits_cache = outmemsys_io_mem_axi_0_aw_bits_cache;
  assign io_mem_axi_0_aw_bits_prot = outmemsys_io_mem_axi_0_aw_bits_prot;
  assign io_mem_axi_0_aw_bits_qos = outmemsys_io_mem_axi_0_aw_bits_qos;
  assign io_mem_axi_0_aw_bits_region = outmemsys_io_mem_axi_0_aw_bits_region;
  assign io_mem_axi_0_aw_bits_id = outmemsys_io_mem_axi_0_aw_bits_id;
  assign io_mem_axi_0_aw_bits_user = outmemsys_io_mem_axi_0_aw_bits_user;
  assign io_mem_axi_0_w_valid = outmemsys_io_mem_axi_0_w_valid;
  assign io_mem_axi_0_w_bits_data = outmemsys_io_mem_axi_0_w_bits_data;
  assign io_mem_axi_0_w_bits_last = outmemsys_io_mem_axi_0_w_bits_last;
  assign io_mem_axi_0_w_bits_id = outmemsys_io_mem_axi_0_w_bits_id;
  assign io_mem_axi_0_w_bits_strb = outmemsys_io_mem_axi_0_w_bits_strb;
  assign io_mem_axi_0_w_bits_user = outmemsys_io_mem_axi_0_w_bits_user;
  assign io_mem_axi_0_b_ready = outmemsys_io_mem_axi_0_b_ready;
  assign io_mem_axi_0_ar_valid = outmemsys_io_mem_axi_0_ar_valid;
  assign io_mem_axi_0_ar_bits_addr = outmemsys_io_mem_axi_0_ar_bits_addr;
  assign io_mem_axi_0_ar_bits_len = outmemsys_io_mem_axi_0_ar_bits_len;
  assign io_mem_axi_0_ar_bits_size = outmemsys_io_mem_axi_0_ar_bits_size;
  assign io_mem_axi_0_ar_bits_burst = outmemsys_io_mem_axi_0_ar_bits_burst;
  assign io_mem_axi_0_ar_bits_lock = outmemsys_io_mem_axi_0_ar_bits_lock;
  assign io_mem_axi_0_ar_bits_cache = outmemsys_io_mem_axi_0_ar_bits_cache;
  assign io_mem_axi_0_ar_bits_prot = outmemsys_io_mem_axi_0_ar_bits_prot;
  assign io_mem_axi_0_ar_bits_qos = outmemsys_io_mem_axi_0_ar_bits_qos;
  assign io_mem_axi_0_ar_bits_region = outmemsys_io_mem_axi_0_ar_bits_region;
  assign io_mem_axi_0_ar_bits_id = outmemsys_io_mem_axi_0_ar_bits_id;
  assign io_mem_axi_0_ar_bits_user = outmemsys_io_mem_axi_0_ar_bits_user;
  assign io_mem_axi_0_r_ready = outmemsys_io_mem_axi_0_r_ready;
  assign io_tiles_cached_0_acquire_ready = outmemsys_io_tiles_cached_0_acquire_ready;
  assign io_tiles_cached_0_probe_valid = outmemsys_io_tiles_cached_0_probe_valid;
  assign io_tiles_cached_0_probe_bits_addr_block = outmemsys_io_tiles_cached_0_probe_bits_addr_block;
  assign io_tiles_cached_0_probe_bits_p_type = outmemsys_io_tiles_cached_0_probe_bits_p_type;
  assign io_tiles_cached_0_release_ready = outmemsys_io_tiles_cached_0_release_ready;
  assign io_tiles_cached_0_grant_valid = outmemsys_io_tiles_cached_0_grant_valid;
  assign io_tiles_cached_0_grant_bits_addr_beat = outmemsys_io_tiles_cached_0_grant_bits_addr_beat;
  assign io_tiles_cached_0_grant_bits_client_xact_id = outmemsys_io_tiles_cached_0_grant_bits_client_xact_id;
  assign io_tiles_cached_0_grant_bits_manager_xact_id = outmemsys_io_tiles_cached_0_grant_bits_manager_xact_id;
  assign io_tiles_cached_0_grant_bits_is_builtin_type = outmemsys_io_tiles_cached_0_grant_bits_is_builtin_type;
  assign io_tiles_cached_0_grant_bits_g_type = outmemsys_io_tiles_cached_0_grant_bits_g_type;
  assign io_tiles_cached_0_grant_bits_data = outmemsys_io_tiles_cached_0_grant_bits_data;
  assign io_tiles_cached_0_grant_bits_manager_id = outmemsys_io_tiles_cached_0_grant_bits_manager_id;
  assign io_tiles_cached_0_finish_ready = outmemsys_io_tiles_cached_0_finish_ready;
  assign io_tiles_uncached_0_acquire_ready = outmemsys_io_tiles_uncached_0_acquire_ready;
  assign io_tiles_uncached_0_grant_valid = outmemsys_io_tiles_uncached_0_grant_valid;
  assign io_tiles_uncached_0_grant_bits_addr_beat = outmemsys_io_tiles_uncached_0_grant_bits_addr_beat;
  assign io_tiles_uncached_0_grant_bits_client_xact_id = outmemsys_io_tiles_uncached_0_grant_bits_client_xact_id;
  assign io_tiles_uncached_0_grant_bits_manager_xact_id = outmemsys_io_tiles_uncached_0_grant_bits_manager_xact_id;
  assign io_tiles_uncached_0_grant_bits_is_builtin_type = outmemsys_io_tiles_uncached_0_grant_bits_is_builtin_type;
  assign io_tiles_uncached_0_grant_bits_g_type = outmemsys_io_tiles_uncached_0_grant_bits_g_type;
  assign io_tiles_uncached_0_grant_bits_data = outmemsys_io_tiles_uncached_0_grant_bits_data;
  assign io_prci_0_reset = reset;
  assign io_prci_0_id = PRCI_1_io_tiles_0_id;
  assign io_prci_0_interrupts_meip = PRCI_1_io_tiles_0_interrupts_meip;
  assign io_prci_0_interrupts_seip = PRCI_1_io_tiles_0_interrupts_seip;
  assign io_prci_0_interrupts_debug = PRCI_1_io_tiles_0_interrupts_debug;
  assign io_prci_0_interrupts_mtip = PRCI_1_io_tiles_0_interrupts_mtip;
  assign io_prci_0_interrupts_msip = PRCI_1_io_tiles_0_interrupts_msip;
  assign io_mmio_axi_0_aw_valid = Queue_19_1_io_deq_valid;
  assign io_mmio_axi_0_aw_bits_addr = Queue_19_1_io_deq_bits_addr;
  assign io_mmio_axi_0_aw_bits_len = Queue_19_1_io_deq_bits_len;
  assign io_mmio_axi_0_aw_bits_size = Queue_19_1_io_deq_bits_size;
  assign io_mmio_axi_0_aw_bits_burst = Queue_19_1_io_deq_bits_burst;
  assign io_mmio_axi_0_aw_bits_lock = Queue_19_1_io_deq_bits_lock;
  assign io_mmio_axi_0_aw_bits_cache = Queue_19_1_io_deq_bits_cache;
  assign io_mmio_axi_0_aw_bits_prot = Queue_19_1_io_deq_bits_prot;
  assign io_mmio_axi_0_aw_bits_qos = Queue_19_1_io_deq_bits_qos;
  assign io_mmio_axi_0_aw_bits_region = Queue_19_1_io_deq_bits_region;
  assign io_mmio_axi_0_aw_bits_id = Queue_19_1_io_deq_bits_id;
  assign io_mmio_axi_0_aw_bits_user = Queue_19_1_io_deq_bits_user;
  assign io_mmio_axi_0_w_valid = Queue_20_1_io_deq_valid;
  assign io_mmio_axi_0_w_bits_data = Queue_20_1_io_deq_bits_data;
  assign io_mmio_axi_0_w_bits_last = Queue_20_1_io_deq_bits_last;
  assign io_mmio_axi_0_w_bits_id = Queue_20_1_io_deq_bits_id;
  assign io_mmio_axi_0_w_bits_strb = Queue_20_1_io_deq_bits_strb;
  assign io_mmio_axi_0_w_bits_user = Queue_20_1_io_deq_bits_user;
  assign io_mmio_axi_0_b_ready = Queue_22_1_io_enq_ready;
  assign io_mmio_axi_0_ar_valid = Queue_18_1_io_deq_valid;
  assign io_mmio_axi_0_ar_bits_addr = Queue_18_1_io_deq_bits_addr;
  assign io_mmio_axi_0_ar_bits_len = Queue_18_1_io_deq_bits_len;
  assign io_mmio_axi_0_ar_bits_size = Queue_18_1_io_deq_bits_size;
  assign io_mmio_axi_0_ar_bits_burst = Queue_18_1_io_deq_bits_burst;
  assign io_mmio_axi_0_ar_bits_lock = Queue_18_1_io_deq_bits_lock;
  assign io_mmio_axi_0_ar_bits_cache = Queue_18_1_io_deq_bits_cache;
  assign io_mmio_axi_0_ar_bits_prot = Queue_18_1_io_deq_bits_prot;
  assign io_mmio_axi_0_ar_bits_qos = Queue_18_1_io_deq_bits_qos;
  assign io_mmio_axi_0_ar_bits_region = Queue_18_1_io_deq_bits_region;
  assign io_mmio_axi_0_ar_bits_id = Queue_18_1_io_deq_bits_id;
  assign io_mmio_axi_0_ar_bits_user = Queue_18_1_io_deq_bits_user;
  assign io_mmio_axi_0_r_ready = Queue_21_1_io_enq_ready;
  assign io_debugBus_req_ready = DebugModule_1_io_db_req_ready;
  assign io_debugBus_resp_valid = DebugModule_1_io_db_resp_valid;
  assign io_debugBus_resp_bits_resp = DebugModule_1_io_db_resp_bits_resp;
  assign io_debugBus_resp_bits_data = DebugModule_1_io_db_resp_bits_data;
  assign outmemsys_clk = clk;
  assign outmemsys_reset = reset;
  assign outmemsys_io_tiles_cached_0_acquire_valid = io_tiles_cached_0_acquire_valid;
  assign outmemsys_io_tiles_cached_0_acquire_bits_addr_block = io_tiles_cached_0_acquire_bits_addr_block;
  assign outmemsys_io_tiles_cached_0_acquire_bits_client_xact_id = io_tiles_cached_0_acquire_bits_client_xact_id;
  assign outmemsys_io_tiles_cached_0_acquire_bits_addr_beat = io_tiles_cached_0_acquire_bits_addr_beat;
  assign outmemsys_io_tiles_cached_0_acquire_bits_is_builtin_type = io_tiles_cached_0_acquire_bits_is_builtin_type;
  assign outmemsys_io_tiles_cached_0_acquire_bits_a_type = io_tiles_cached_0_acquire_bits_a_type;
  assign outmemsys_io_tiles_cached_0_acquire_bits_union = io_tiles_cached_0_acquire_bits_union;
  assign outmemsys_io_tiles_cached_0_acquire_bits_data = io_tiles_cached_0_acquire_bits_data;
  assign outmemsys_io_tiles_cached_0_probe_ready = io_tiles_cached_0_probe_ready;
  assign outmemsys_io_tiles_cached_0_release_valid = io_tiles_cached_0_release_valid;
  assign outmemsys_io_tiles_cached_0_release_bits_addr_beat = io_tiles_cached_0_release_bits_addr_beat;
  assign outmemsys_io_tiles_cached_0_release_bits_addr_block = io_tiles_cached_0_release_bits_addr_block;
  assign outmemsys_io_tiles_cached_0_release_bits_client_xact_id = io_tiles_cached_0_release_bits_client_xact_id;
  assign outmemsys_io_tiles_cached_0_release_bits_voluntary = io_tiles_cached_0_release_bits_voluntary;
  assign outmemsys_io_tiles_cached_0_release_bits_r_type = io_tiles_cached_0_release_bits_r_type;
  assign outmemsys_io_tiles_cached_0_release_bits_data = io_tiles_cached_0_release_bits_data;
  assign outmemsys_io_tiles_cached_0_grant_ready = io_tiles_cached_0_grant_ready;
  assign outmemsys_io_tiles_cached_0_finish_valid = io_tiles_cached_0_finish_valid;
  assign outmemsys_io_tiles_cached_0_finish_bits_manager_xact_id = io_tiles_cached_0_finish_bits_manager_xact_id;
  assign outmemsys_io_tiles_cached_0_finish_bits_manager_id = io_tiles_cached_0_finish_bits_manager_id;
  assign outmemsys_io_tiles_uncached_0_acquire_valid = io_tiles_uncached_0_acquire_valid;
  assign outmemsys_io_tiles_uncached_0_acquire_bits_addr_block = io_tiles_uncached_0_acquire_bits_addr_block;
  assign outmemsys_io_tiles_uncached_0_acquire_bits_client_xact_id = io_tiles_uncached_0_acquire_bits_client_xact_id;
  assign outmemsys_io_tiles_uncached_0_acquire_bits_addr_beat = io_tiles_uncached_0_acquire_bits_addr_beat;
  assign outmemsys_io_tiles_uncached_0_acquire_bits_is_builtin_type = io_tiles_uncached_0_acquire_bits_is_builtin_type;
  assign outmemsys_io_tiles_uncached_0_acquire_bits_a_type = io_tiles_uncached_0_acquire_bits_a_type;
  assign outmemsys_io_tiles_uncached_0_acquire_bits_union = io_tiles_uncached_0_acquire_bits_union;
  assign outmemsys_io_tiles_uncached_0_acquire_bits_data = io_tiles_uncached_0_acquire_bits_data;
  assign outmemsys_io_tiles_uncached_0_grant_ready = io_tiles_uncached_0_grant_ready;
  assign outmemsys_io_incoherent_0 = 1'h0;
  assign outmemsys_io_mem_axi_0_aw_ready = io_mem_axi_0_aw_ready;
  assign outmemsys_io_mem_axi_0_w_ready = io_mem_axi_0_w_ready;
  assign outmemsys_io_mem_axi_0_b_valid = io_mem_axi_0_b_valid;
  assign outmemsys_io_mem_axi_0_b_bits_resp = io_mem_axi_0_b_bits_resp;
  assign outmemsys_io_mem_axi_0_b_bits_id = io_mem_axi_0_b_bits_id;
  assign outmemsys_io_mem_axi_0_b_bits_user = io_mem_axi_0_b_bits_user;
  assign outmemsys_io_mem_axi_0_ar_ready = io_mem_axi_0_ar_ready;
  assign outmemsys_io_mem_axi_0_r_valid = io_mem_axi_0_r_valid;
  assign outmemsys_io_mem_axi_0_r_bits_resp = io_mem_axi_0_r_bits_resp;
  assign outmemsys_io_mem_axi_0_r_bits_data = io_mem_axi_0_r_bits_data;
  assign outmemsys_io_mem_axi_0_r_bits_last = io_mem_axi_0_r_bits_last;
  assign outmemsys_io_mem_axi_0_r_bits_id = io_mem_axi_0_r_bits_id;
  assign outmemsys_io_mem_axi_0_r_bits_user = io_mem_axi_0_r_bits_user;
  assign outmemsys_io_mmio_acquire_ready = TileLinkRecursiveInterconnect_2_io_in_0_acquire_ready;
  assign outmemsys_io_mmio_grant_valid = TileLinkRecursiveInterconnect_2_io_in_0_grant_valid;
  assign outmemsys_io_mmio_grant_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_addr_beat;
  assign outmemsys_io_mmio_grant_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_client_xact_id;
  assign outmemsys_io_mmio_grant_bits_manager_xact_id = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_manager_xact_id;
  assign outmemsys_io_mmio_grant_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_is_builtin_type;
  assign outmemsys_io_mmio_grant_bits_g_type = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_g_type;
  assign outmemsys_io_mmio_grant_bits_data = TileLinkRecursiveInterconnect_2_io_in_0_grant_bits_data;
  assign TileLinkRecursiveInterconnect_2_clk = clk;
  assign TileLinkRecursiveInterconnect_2_reset = reset;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_valid = outmemsys_io_mmio_acquire_valid;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_block = outmemsys_io_mmio_acquire_bits_addr_block;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_client_xact_id = outmemsys_io_mmio_acquire_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_addr_beat = outmemsys_io_mmio_acquire_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_is_builtin_type = outmemsys_io_mmio_acquire_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_a_type = outmemsys_io_mmio_acquire_bits_a_type;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_union = outmemsys_io_mmio_acquire_bits_union;
  assign TileLinkRecursiveInterconnect_2_io_in_0_acquire_bits_data = outmemsys_io_mmio_acquire_bits_data;
  assign TileLinkRecursiveInterconnect_2_io_in_0_grant_ready = outmemsys_io_mmio_grant_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_0_acquire_ready = DebugModule_1_io_tl_acquire_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_valid = DebugModule_1_io_tl_grant_valid;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_addr_beat = DebugModule_1_io_tl_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_client_xact_id = DebugModule_1_io_tl_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_manager_xact_id = DebugModule_1_io_tl_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_is_builtin_type = DebugModule_1_io_tl_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_g_type = DebugModule_1_io_tl_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_2_io_out_0_grant_bits_data = DebugModule_1_io_tl_grant_bits_data;
  assign TileLinkRecursiveInterconnect_2_io_out_1_acquire_ready = ROMSlave_1_io_acquire_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_valid = ROMSlave_1_io_grant_valid;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_addr_beat = ROMSlave_1_io_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_client_xact_id = ROMSlave_1_io_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_manager_xact_id = ROMSlave_1_io_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_is_builtin_type = ROMSlave_1_io_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_g_type = ROMSlave_1_io_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_2_io_out_1_grant_bits_data = ROMSlave_1_io_grant_bits_data;
  assign TileLinkRecursiveInterconnect_2_io_out_2_acquire_ready = PLIC_1_io_tl_acquire_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_valid = PLIC_1_io_tl_grant_valid;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_addr_beat = PLIC_1_io_tl_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_client_xact_id = PLIC_1_io_tl_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_manager_xact_id = PLIC_1_io_tl_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_is_builtin_type = PLIC_1_io_tl_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_g_type = PLIC_1_io_tl_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_2_io_out_2_grant_bits_data = PLIC_1_io_tl_grant_bits_data;
  assign TileLinkRecursiveInterconnect_2_io_out_3_acquire_ready = PRCI_1_io_tl_acquire_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_valid = PRCI_1_io_tl_grant_valid;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_addr_beat = PRCI_1_io_tl_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_client_xact_id = PRCI_1_io_tl_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_manager_xact_id = PRCI_1_io_tl_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_is_builtin_type = PRCI_1_io_tl_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_g_type = PRCI_1_io_tl_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_2_io_out_3_grant_bits_data = PRCI_1_io_tl_grant_bits_data;
  assign TileLinkRecursiveInterconnect_2_io_out_4_acquire_ready = NastiIOTileLinkIOConverter_1_1_io_tl_acquire_ready;
  assign TileLinkRecursiveInterconnect_2_io_out_4_grant_valid = NastiIOTileLinkIOConverter_1_1_io_tl_grant_valid;
  assign TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_addr_beat = NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_client_xact_id = NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_manager_xact_id = NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_is_builtin_type = NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_g_type = NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_2_io_out_4_grant_bits_data = NastiIOTileLinkIOConverter_1_1_io_tl_grant_bits_data;
  assign PLIC_1_clk = clk;
  assign PLIC_1_reset = reset;
  assign PLIC_1_io_devices_0_valid = LevelGateway_31_io_plic_valid;
  assign PLIC_1_io_devices_1_valid = LevelGateway_1_1_io_plic_valid;
  assign PLIC_1_io_devices_2_valid = LevelGateway_2_1_io_plic_valid;
  assign PLIC_1_io_devices_3_valid = LevelGateway_3_1_io_plic_valid;
  assign PLIC_1_io_devices_4_valid = LevelGateway_4_1_io_plic_valid;
  assign PLIC_1_io_devices_5_valid = LevelGateway_5_1_io_plic_valid;
  assign PLIC_1_io_devices_6_valid = LevelGateway_6_1_io_plic_valid;
  assign PLIC_1_io_devices_7_valid = LevelGateway_7_1_io_plic_valid;
  assign PLIC_1_io_devices_8_valid = LevelGateway_8_1_io_plic_valid;
  assign PLIC_1_io_devices_9_valid = LevelGateway_9_1_io_plic_valid;
  assign PLIC_1_io_devices_10_valid = LevelGateway_10_1_io_plic_valid;
  assign PLIC_1_io_devices_11_valid = LevelGateway_11_1_io_plic_valid;
  assign PLIC_1_io_devices_12_valid = LevelGateway_12_1_io_plic_valid;
  assign PLIC_1_io_devices_13_valid = LevelGateway_13_1_io_plic_valid;
  assign PLIC_1_io_devices_14_valid = LevelGateway_14_1_io_plic_valid;
  assign PLIC_1_io_devices_15_valid = LevelGateway_15_1_io_plic_valid;
  assign PLIC_1_io_devices_16_valid = LevelGateway_16_1_io_plic_valid;
  assign PLIC_1_io_devices_17_valid = LevelGateway_17_1_io_plic_valid;
  assign PLIC_1_io_devices_18_valid = LevelGateway_18_1_io_plic_valid;
  assign PLIC_1_io_devices_19_valid = LevelGateway_19_1_io_plic_valid;
  assign PLIC_1_io_devices_20_valid = LevelGateway_20_1_io_plic_valid;
  assign PLIC_1_io_devices_21_valid = LevelGateway_21_1_io_plic_valid;
  assign PLIC_1_io_devices_22_valid = LevelGateway_22_1_io_plic_valid;
  assign PLIC_1_io_devices_23_valid = LevelGateway_23_1_io_plic_valid;
  assign PLIC_1_io_devices_24_valid = LevelGateway_24_1_io_plic_valid;
  assign PLIC_1_io_devices_25_valid = LevelGateway_25_1_io_plic_valid;
  assign PLIC_1_io_devices_26_valid = LevelGateway_26_1_io_plic_valid;
  assign PLIC_1_io_devices_27_valid = LevelGateway_27_1_io_plic_valid;
  assign PLIC_1_io_devices_28_valid = LevelGateway_28_1_io_plic_valid;
  assign PLIC_1_io_devices_29_valid = LevelGateway_29_1_io_plic_valid;
  assign PLIC_1_io_devices_30_valid = LevelGateway_30_1_io_plic_valid;
  assign PLIC_1_io_tl_acquire_valid = TileLinkRecursiveInterconnect_2_io_out_2_acquire_valid;
  assign PLIC_1_io_tl_acquire_bits_addr_block = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_block;
  assign PLIC_1_io_tl_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_client_xact_id;
  assign PLIC_1_io_tl_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_addr_beat;
  assign PLIC_1_io_tl_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_is_builtin_type;
  assign PLIC_1_io_tl_acquire_bits_a_type = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_a_type;
  assign PLIC_1_io_tl_acquire_bits_union = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_union;
  assign PLIC_1_io_tl_acquire_bits_data = TileLinkRecursiveInterconnect_2_io_out_2_acquire_bits_data;
  assign PLIC_1_io_tl_grant_ready = TileLinkRecursiveInterconnect_2_io_out_2_grant_ready;
  assign LevelGateway_31_clk = clk;
  assign LevelGateway_31_reset = reset;
  assign LevelGateway_31_io_interrupt = io_interrupts_0;
  assign LevelGateway_31_io_plic_ready = PLIC_1_io_devices_0_ready;
  assign LevelGateway_31_io_plic_complete = PLIC_1_io_devices_0_complete;
  assign LevelGateway_1_1_clk = clk;
  assign LevelGateway_1_1_reset = reset;
  assign LevelGateway_1_1_io_interrupt = io_interrupts_1;
  assign LevelGateway_1_1_io_plic_ready = PLIC_1_io_devices_1_ready;
  assign LevelGateway_1_1_io_plic_complete = PLIC_1_io_devices_1_complete;
  assign LevelGateway_2_1_clk = clk;
  assign LevelGateway_2_1_reset = reset;
  assign LevelGateway_2_1_io_interrupt = io_interrupts_2;
  assign LevelGateway_2_1_io_plic_ready = PLIC_1_io_devices_2_ready;
  assign LevelGateway_2_1_io_plic_complete = PLIC_1_io_devices_2_complete;
  assign LevelGateway_3_1_clk = clk;
  assign LevelGateway_3_1_reset = reset;
  assign LevelGateway_3_1_io_interrupt = io_interrupts_3;
  assign LevelGateway_3_1_io_plic_ready = PLIC_1_io_devices_3_ready;
  assign LevelGateway_3_1_io_plic_complete = PLIC_1_io_devices_3_complete;
  assign LevelGateway_4_1_clk = clk;
  assign LevelGateway_4_1_reset = reset;
  assign LevelGateway_4_1_io_interrupt = io_interrupts_4;
  assign LevelGateway_4_1_io_plic_ready = PLIC_1_io_devices_4_ready;
  assign LevelGateway_4_1_io_plic_complete = PLIC_1_io_devices_4_complete;
  assign LevelGateway_5_1_clk = clk;
  assign LevelGateway_5_1_reset = reset;
  assign LevelGateway_5_1_io_interrupt = io_interrupts_5;
  assign LevelGateway_5_1_io_plic_ready = PLIC_1_io_devices_5_ready;
  assign LevelGateway_5_1_io_plic_complete = PLIC_1_io_devices_5_complete;
  assign LevelGateway_6_1_clk = clk;
  assign LevelGateway_6_1_reset = reset;
  assign LevelGateway_6_1_io_interrupt = io_interrupts_6;
  assign LevelGateway_6_1_io_plic_ready = PLIC_1_io_devices_6_ready;
  assign LevelGateway_6_1_io_plic_complete = PLIC_1_io_devices_6_complete;
  assign LevelGateway_7_1_clk = clk;
  assign LevelGateway_7_1_reset = reset;
  assign LevelGateway_7_1_io_interrupt = io_interrupts_7;
  assign LevelGateway_7_1_io_plic_ready = PLIC_1_io_devices_7_ready;
  assign LevelGateway_7_1_io_plic_complete = PLIC_1_io_devices_7_complete;
  assign LevelGateway_8_1_clk = clk;
  assign LevelGateway_8_1_reset = reset;
  assign LevelGateway_8_1_io_interrupt = io_interrupts_8;
  assign LevelGateway_8_1_io_plic_ready = PLIC_1_io_devices_8_ready;
  assign LevelGateway_8_1_io_plic_complete = PLIC_1_io_devices_8_complete;
  assign LevelGateway_9_1_clk = clk;
  assign LevelGateway_9_1_reset = reset;
  assign LevelGateway_9_1_io_interrupt = io_interrupts_9;
  assign LevelGateway_9_1_io_plic_ready = PLIC_1_io_devices_9_ready;
  assign LevelGateway_9_1_io_plic_complete = PLIC_1_io_devices_9_complete;
  assign LevelGateway_10_1_clk = clk;
  assign LevelGateway_10_1_reset = reset;
  assign LevelGateway_10_1_io_interrupt = io_interrupts_10;
  assign LevelGateway_10_1_io_plic_ready = PLIC_1_io_devices_10_ready;
  assign LevelGateway_10_1_io_plic_complete = PLIC_1_io_devices_10_complete;
  assign LevelGateway_11_1_clk = clk;
  assign LevelGateway_11_1_reset = reset;
  assign LevelGateway_11_1_io_interrupt = io_interrupts_11;
  assign LevelGateway_11_1_io_plic_ready = PLIC_1_io_devices_11_ready;
  assign LevelGateway_11_1_io_plic_complete = PLIC_1_io_devices_11_complete;
  assign LevelGateway_12_1_clk = clk;
  assign LevelGateway_12_1_reset = reset;
  assign LevelGateway_12_1_io_interrupt = io_interrupts_12;
  assign LevelGateway_12_1_io_plic_ready = PLIC_1_io_devices_12_ready;
  assign LevelGateway_12_1_io_plic_complete = PLIC_1_io_devices_12_complete;
  assign LevelGateway_13_1_clk = clk;
  assign LevelGateway_13_1_reset = reset;
  assign LevelGateway_13_1_io_interrupt = io_interrupts_13;
  assign LevelGateway_13_1_io_plic_ready = PLIC_1_io_devices_13_ready;
  assign LevelGateway_13_1_io_plic_complete = PLIC_1_io_devices_13_complete;
  assign LevelGateway_14_1_clk = clk;
  assign LevelGateway_14_1_reset = reset;
  assign LevelGateway_14_1_io_interrupt = io_interrupts_14;
  assign LevelGateway_14_1_io_plic_ready = PLIC_1_io_devices_14_ready;
  assign LevelGateway_14_1_io_plic_complete = PLIC_1_io_devices_14_complete;
  assign LevelGateway_15_1_clk = clk;
  assign LevelGateway_15_1_reset = reset;
  assign LevelGateway_15_1_io_interrupt = io_interrupts_15;
  assign LevelGateway_15_1_io_plic_ready = PLIC_1_io_devices_15_ready;
  assign LevelGateway_15_1_io_plic_complete = PLIC_1_io_devices_15_complete;
  assign LevelGateway_16_1_clk = clk;
  assign LevelGateway_16_1_reset = reset;
  assign LevelGateway_16_1_io_interrupt = io_interrupts_16;
  assign LevelGateway_16_1_io_plic_ready = PLIC_1_io_devices_16_ready;
  assign LevelGateway_16_1_io_plic_complete = PLIC_1_io_devices_16_complete;
  assign LevelGateway_17_1_clk = clk;
  assign LevelGateway_17_1_reset = reset;
  assign LevelGateway_17_1_io_interrupt = io_interrupts_17;
  assign LevelGateway_17_1_io_plic_ready = PLIC_1_io_devices_17_ready;
  assign LevelGateway_17_1_io_plic_complete = PLIC_1_io_devices_17_complete;
  assign LevelGateway_18_1_clk = clk;
  assign LevelGateway_18_1_reset = reset;
  assign LevelGateway_18_1_io_interrupt = io_interrupts_18;
  assign LevelGateway_18_1_io_plic_ready = PLIC_1_io_devices_18_ready;
  assign LevelGateway_18_1_io_plic_complete = PLIC_1_io_devices_18_complete;
  assign LevelGateway_19_1_clk = clk;
  assign LevelGateway_19_1_reset = reset;
  assign LevelGateway_19_1_io_interrupt = io_interrupts_19;
  assign LevelGateway_19_1_io_plic_ready = PLIC_1_io_devices_19_ready;
  assign LevelGateway_19_1_io_plic_complete = PLIC_1_io_devices_19_complete;
  assign LevelGateway_20_1_clk = clk;
  assign LevelGateway_20_1_reset = reset;
  assign LevelGateway_20_1_io_interrupt = io_interrupts_20;
  assign LevelGateway_20_1_io_plic_ready = PLIC_1_io_devices_20_ready;
  assign LevelGateway_20_1_io_plic_complete = PLIC_1_io_devices_20_complete;
  assign LevelGateway_21_1_clk = clk;
  assign LevelGateway_21_1_reset = reset;
  assign LevelGateway_21_1_io_interrupt = io_interrupts_21;
  assign LevelGateway_21_1_io_plic_ready = PLIC_1_io_devices_21_ready;
  assign LevelGateway_21_1_io_plic_complete = PLIC_1_io_devices_21_complete;
  assign LevelGateway_22_1_clk = clk;
  assign LevelGateway_22_1_reset = reset;
  assign LevelGateway_22_1_io_interrupt = io_interrupts_22;
  assign LevelGateway_22_1_io_plic_ready = PLIC_1_io_devices_22_ready;
  assign LevelGateway_22_1_io_plic_complete = PLIC_1_io_devices_22_complete;
  assign LevelGateway_23_1_clk = clk;
  assign LevelGateway_23_1_reset = reset;
  assign LevelGateway_23_1_io_interrupt = io_interrupts_23;
  assign LevelGateway_23_1_io_plic_ready = PLIC_1_io_devices_23_ready;
  assign LevelGateway_23_1_io_plic_complete = PLIC_1_io_devices_23_complete;
  assign LevelGateway_24_1_clk = clk;
  assign LevelGateway_24_1_reset = reset;
  assign LevelGateway_24_1_io_interrupt = io_interrupts_24;
  assign LevelGateway_24_1_io_plic_ready = PLIC_1_io_devices_24_ready;
  assign LevelGateway_24_1_io_plic_complete = PLIC_1_io_devices_24_complete;
  assign LevelGateway_25_1_clk = clk;
  assign LevelGateway_25_1_reset = reset;
  assign LevelGateway_25_1_io_interrupt = io_interrupts_25;
  assign LevelGateway_25_1_io_plic_ready = PLIC_1_io_devices_25_ready;
  assign LevelGateway_25_1_io_plic_complete = PLIC_1_io_devices_25_complete;
  assign LevelGateway_26_1_clk = clk;
  assign LevelGateway_26_1_reset = reset;
  assign LevelGateway_26_1_io_interrupt = io_interrupts_26;
  assign LevelGateway_26_1_io_plic_ready = PLIC_1_io_devices_26_ready;
  assign LevelGateway_26_1_io_plic_complete = PLIC_1_io_devices_26_complete;
  assign LevelGateway_27_1_clk = clk;
  assign LevelGateway_27_1_reset = reset;
  assign LevelGateway_27_1_io_interrupt = io_interrupts_27;
  assign LevelGateway_27_1_io_plic_ready = PLIC_1_io_devices_27_ready;
  assign LevelGateway_27_1_io_plic_complete = PLIC_1_io_devices_27_complete;
  assign LevelGateway_28_1_clk = clk;
  assign LevelGateway_28_1_reset = reset;
  assign LevelGateway_28_1_io_interrupt = io_interrupts_28;
  assign LevelGateway_28_1_io_plic_ready = PLIC_1_io_devices_28_ready;
  assign LevelGateway_28_1_io_plic_complete = PLIC_1_io_devices_28_complete;
  assign LevelGateway_29_1_clk = clk;
  assign LevelGateway_29_1_reset = reset;
  assign LevelGateway_29_1_io_interrupt = io_interrupts_29;
  assign LevelGateway_29_1_io_plic_ready = PLIC_1_io_devices_29_ready;
  assign LevelGateway_29_1_io_plic_complete = PLIC_1_io_devices_29_complete;
  assign LevelGateway_30_1_clk = clk;
  assign LevelGateway_30_1_reset = reset;
  assign LevelGateway_30_1_io_interrupt = io_interrupts_30;
  assign LevelGateway_30_1_io_plic_ready = PLIC_1_io_devices_30_ready;
  assign LevelGateway_30_1_io_plic_complete = PLIC_1_io_devices_30_complete;
  assign DebugModule_1_clk = clk;
  assign DebugModule_1_reset = reset;
  assign DebugModule_1_io_db_req_valid = io_debugBus_req_valid;
  assign DebugModule_1_io_db_req_bits_addr = io_debugBus_req_bits_addr;
  assign DebugModule_1_io_db_req_bits_op = io_debugBus_req_bits_op;
  assign DebugModule_1_io_db_req_bits_data = io_debugBus_req_bits_data;
  assign DebugModule_1_io_db_resp_ready = io_debugBus_resp_ready;
  assign DebugModule_1_io_tl_acquire_valid = TileLinkRecursiveInterconnect_2_io_out_0_acquire_valid;
  assign DebugModule_1_io_tl_acquire_bits_addr_block = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_block;
  assign DebugModule_1_io_tl_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_client_xact_id;
  assign DebugModule_1_io_tl_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_addr_beat;
  assign DebugModule_1_io_tl_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_is_builtin_type;
  assign DebugModule_1_io_tl_acquire_bits_a_type = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_a_type;
  assign DebugModule_1_io_tl_acquire_bits_union = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_union;
  assign DebugModule_1_io_tl_acquire_bits_data = TileLinkRecursiveInterconnect_2_io_out_0_acquire_bits_data;
  assign DebugModule_1_io_tl_grant_ready = TileLinkRecursiveInterconnect_2_io_out_0_grant_ready;
  assign PRCI_1_clk = clk;
  assign PRCI_1_reset = reset;
  assign PRCI_1_io_interrupts_0_meip = PLIC_1_io_harts_0;
  assign PRCI_1_io_interrupts_0_seip = GEN_1;
  assign PRCI_1_io_interrupts_0_debug = DebugModule_1_io_debugInterrupts_0;
  assign PRCI_1_io_tl_acquire_valid = TileLinkRecursiveInterconnect_2_io_out_3_acquire_valid;
  assign PRCI_1_io_tl_acquire_bits_addr_block = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_block;
  assign PRCI_1_io_tl_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_client_xact_id;
  assign PRCI_1_io_tl_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_addr_beat;
  assign PRCI_1_io_tl_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_is_builtin_type;
  assign PRCI_1_io_tl_acquire_bits_a_type = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_a_type;
  assign PRCI_1_io_tl_acquire_bits_union = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_union;
  assign PRCI_1_io_tl_acquire_bits_data = TileLinkRecursiveInterconnect_2_io_out_3_acquire_bits_data;
  assign PRCI_1_io_tl_grant_ready = TileLinkRecursiveInterconnect_2_io_out_3_grant_ready;
  assign PRCI_1_io_rtcTick = T_10391;
  assign T_10391 = T_10389 == 7'h63;
  assign T_10393 = T_10389 + 7'h1;
  assign T_10394 = T_10393[6:0];
  assign GEN_0 = T_10391 ? 7'h0 : T_10394;
  assign ROMSlave_1_clk = clk;
  assign ROMSlave_1_reset = reset;
  assign ROMSlave_1_io_acquire_valid = TileLinkRecursiveInterconnect_2_io_out_1_acquire_valid;
  assign ROMSlave_1_io_acquire_bits_addr_block = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_block;
  assign ROMSlave_1_io_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_client_xact_id;
  assign ROMSlave_1_io_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_addr_beat;
  assign ROMSlave_1_io_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_is_builtin_type;
  assign ROMSlave_1_io_acquire_bits_a_type = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_a_type;
  assign ROMSlave_1_io_acquire_bits_union = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_union;
  assign ROMSlave_1_io_acquire_bits_data = TileLinkRecursiveInterconnect_2_io_out_1_acquire_bits_data;
  assign ROMSlave_1_io_grant_ready = TileLinkRecursiveInterconnect_2_io_out_1_grant_ready;
  assign NastiIOTileLinkIOConverter_1_1_clk = clk;
  assign NastiIOTileLinkIOConverter_1_1_reset = reset;
  assign NastiIOTileLinkIOConverter_1_1_io_tl_acquire_valid = TileLinkRecursiveInterconnect_2_io_out_4_acquire_valid;
  assign NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_addr_block = TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_addr_block;
  assign NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_client_xact_id;
  assign NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_addr_beat;
  assign NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_is_builtin_type;
  assign NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_a_type = TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_a_type;
  assign NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_union = TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_union;
  assign NastiIOTileLinkIOConverter_1_1_io_tl_acquire_bits_data = TileLinkRecursiveInterconnect_2_io_out_4_acquire_bits_data;
  assign NastiIOTileLinkIOConverter_1_1_io_tl_grant_ready = TileLinkRecursiveInterconnect_2_io_out_4_grant_ready;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_aw_ready = Queue_19_1_io_enq_ready;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_w_ready = Queue_20_1_io_enq_ready;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_b_valid = Queue_22_1_io_deq_valid;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_b_bits_resp = Queue_22_1_io_deq_bits_resp;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_b_bits_id = Queue_22_1_io_deq_bits_id;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_b_bits_user = Queue_22_1_io_deq_bits_user;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_ar_ready = Queue_18_1_io_enq_ready;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_r_valid = Queue_21_1_io_deq_valid;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_resp = Queue_21_1_io_deq_bits_resp;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_data = Queue_21_1_io_deq_bits_data;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_last = Queue_21_1_io_deq_bits_last;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_id = Queue_21_1_io_deq_bits_id;
  assign NastiIOTileLinkIOConverter_1_1_io_nasti_r_bits_user = Queue_21_1_io_deq_bits_user;
  assign Queue_18_1_clk = clk;
  assign Queue_18_1_reset = reset;
  assign Queue_18_1_io_enq_valid = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_valid;
  assign Queue_18_1_io_enq_bits_addr = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_addr;
  assign Queue_18_1_io_enq_bits_len = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_len;
  assign Queue_18_1_io_enq_bits_size = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_size;
  assign Queue_18_1_io_enq_bits_burst = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_burst;
  assign Queue_18_1_io_enq_bits_lock = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_lock;
  assign Queue_18_1_io_enq_bits_cache = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_cache;
  assign Queue_18_1_io_enq_bits_prot = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_prot;
  assign Queue_18_1_io_enq_bits_qos = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_qos;
  assign Queue_18_1_io_enq_bits_region = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_region;
  assign Queue_18_1_io_enq_bits_id = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_id;
  assign Queue_18_1_io_enq_bits_user = NastiIOTileLinkIOConverter_1_1_io_nasti_ar_bits_user;
  assign Queue_18_1_io_deq_ready = io_mmio_axi_0_ar_ready;
  assign Queue_19_1_clk = clk;
  assign Queue_19_1_reset = reset;
  assign Queue_19_1_io_enq_valid = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_valid;
  assign Queue_19_1_io_enq_bits_addr = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_addr;
  assign Queue_19_1_io_enq_bits_len = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_len;
  assign Queue_19_1_io_enq_bits_size = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_size;
  assign Queue_19_1_io_enq_bits_burst = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_burst;
  assign Queue_19_1_io_enq_bits_lock = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_lock;
  assign Queue_19_1_io_enq_bits_cache = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_cache;
  assign Queue_19_1_io_enq_bits_prot = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_prot;
  assign Queue_19_1_io_enq_bits_qos = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_qos;
  assign Queue_19_1_io_enq_bits_region = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_region;
  assign Queue_19_1_io_enq_bits_id = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_id;
  assign Queue_19_1_io_enq_bits_user = NastiIOTileLinkIOConverter_1_1_io_nasti_aw_bits_user;
  assign Queue_19_1_io_deq_ready = io_mmio_axi_0_aw_ready;
  assign Queue_20_1_clk = clk;
  assign Queue_20_1_reset = reset;
  assign Queue_20_1_io_enq_valid = NastiIOTileLinkIOConverter_1_1_io_nasti_w_valid;
  assign Queue_20_1_io_enq_bits_data = NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_data;
  assign Queue_20_1_io_enq_bits_last = NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_last;
  assign Queue_20_1_io_enq_bits_id = NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_id;
  assign Queue_20_1_io_enq_bits_strb = NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_strb;
  assign Queue_20_1_io_enq_bits_user = NastiIOTileLinkIOConverter_1_1_io_nasti_w_bits_user;
  assign Queue_20_1_io_deq_ready = io_mmio_axi_0_w_ready;
  assign Queue_21_1_clk = clk;
  assign Queue_21_1_reset = reset;
  assign Queue_21_1_io_enq_valid = io_mmio_axi_0_r_valid;
  assign Queue_21_1_io_enq_bits_resp = io_mmio_axi_0_r_bits_resp;
  assign Queue_21_1_io_enq_bits_data = io_mmio_axi_0_r_bits_data;
  assign Queue_21_1_io_enq_bits_last = io_mmio_axi_0_r_bits_last;
  assign Queue_21_1_io_enq_bits_id = io_mmio_axi_0_r_bits_id;
  assign Queue_21_1_io_enq_bits_user = io_mmio_axi_0_r_bits_user;
  assign Queue_21_1_io_deq_ready = NastiIOTileLinkIOConverter_1_1_io_nasti_r_ready;
  assign Queue_22_1_clk = clk;
  assign Queue_22_1_reset = reset;
  assign Queue_22_1_io_enq_valid = io_mmio_axi_0_b_valid;
  assign Queue_22_1_io_enq_bits_resp = io_mmio_axi_0_b_bits_resp;
  assign Queue_22_1_io_enq_bits_id = io_mmio_axi_0_b_bits_id;
  assign Queue_22_1_io_enq_bits_user = io_mmio_axi_0_b_bits_user;
  assign Queue_22_1_io_deq_ready = NastiIOTileLinkIOConverter_1_1_io_nasti_b_ready;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_2 = {1{$random}};
  T_10389 = GEN_2[6:0];
  `endif
  `ifdef RANDOMIZE
  GEN_3 = {1{$random}};
  GEN_1 = GEN_3[0:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_10389 <= 7'h0;
    end else begin
      if(T_10391) begin
        T_10389 <= 7'h0;
      end else begin
        T_10389 <= T_10394;
      end
    end
  end
endmodule
module Top(
  input   clk,
  input   reset,
  input   io_mem_axi_0_aw_ready,
  output  io_mem_axi_0_aw_valid,
  output [31:0] io_mem_axi_0_aw_bits_addr,
  output [7:0] io_mem_axi_0_aw_bits_len,
  output [2:0] io_mem_axi_0_aw_bits_size,
  output [1:0] io_mem_axi_0_aw_bits_burst,
  output  io_mem_axi_0_aw_bits_lock,
  output [3:0] io_mem_axi_0_aw_bits_cache,
  output [2:0] io_mem_axi_0_aw_bits_prot,
  output [3:0] io_mem_axi_0_aw_bits_qos,
  output [3:0] io_mem_axi_0_aw_bits_region,
  output [4:0] io_mem_axi_0_aw_bits_id,
  output  io_mem_axi_0_aw_bits_user,
  input   io_mem_axi_0_w_ready,
  output  io_mem_axi_0_w_valid,
  output [63:0] io_mem_axi_0_w_bits_data,
  output  io_mem_axi_0_w_bits_last,
  output [4:0] io_mem_axi_0_w_bits_id,
  output [7:0] io_mem_axi_0_w_bits_strb,
  output  io_mem_axi_0_w_bits_user,
  output  io_mem_axi_0_b_ready,
  input   io_mem_axi_0_b_valid,
  input  [1:0] io_mem_axi_0_b_bits_resp,
  input  [4:0] io_mem_axi_0_b_bits_id,
  input   io_mem_axi_0_b_bits_user,
  input   io_mem_axi_0_ar_ready,
  output  io_mem_axi_0_ar_valid,
  output [31:0] io_mem_axi_0_ar_bits_addr,
  output [7:0] io_mem_axi_0_ar_bits_len,
  output [2:0] io_mem_axi_0_ar_bits_size,
  output [1:0] io_mem_axi_0_ar_bits_burst,
  output  io_mem_axi_0_ar_bits_lock,
  output [3:0] io_mem_axi_0_ar_bits_cache,
  output [2:0] io_mem_axi_0_ar_bits_prot,
  output [3:0] io_mem_axi_0_ar_bits_qos,
  output [3:0] io_mem_axi_0_ar_bits_region,
  output [4:0] io_mem_axi_0_ar_bits_id,
  output  io_mem_axi_0_ar_bits_user,
  output  io_mem_axi_0_r_ready,
  input   io_mem_axi_0_r_valid,
  input  [1:0] io_mem_axi_0_r_bits_resp,
  input  [63:0] io_mem_axi_0_r_bits_data,
  input   io_mem_axi_0_r_bits_last,
  input  [4:0] io_mem_axi_0_r_bits_id,
  input   io_mem_axi_0_r_bits_user,
  input   io_interrupts_0,
  input   io_interrupts_1,
  input   io_interrupts_2,
  input   io_interrupts_3,
  input   io_interrupts_4,
  input   io_interrupts_5,
  input   io_interrupts_6,
  input   io_interrupts_7,
  input   io_interrupts_8,
  input   io_interrupts_9,
  input   io_interrupts_10,
  input   io_interrupts_11,
  input   io_interrupts_12,
  input   io_interrupts_13,
  input   io_interrupts_14,
  input   io_interrupts_15,
  input   io_interrupts_16,
  input   io_interrupts_17,
  input   io_interrupts_18,
  input   io_interrupts_19,
  input   io_interrupts_20,
  input   io_interrupts_21,
  input   io_interrupts_22,
  input   io_interrupts_23,
  input   io_interrupts_24,
  input   io_interrupts_25,
  input   io_interrupts_26,
  input   io_interrupts_27,
  input   io_interrupts_28,
  input   io_interrupts_29,
  input   io_interrupts_30,
  input   io_mmio_axi_0_aw_ready,
  output  io_mmio_axi_0_aw_valid,
  output [31:0] io_mmio_axi_0_aw_bits_addr,
  output [7:0] io_mmio_axi_0_aw_bits_len,
  output [2:0] io_mmio_axi_0_aw_bits_size,
  output [1:0] io_mmio_axi_0_aw_bits_burst,
  output  io_mmio_axi_0_aw_bits_lock,
  output [3:0] io_mmio_axi_0_aw_bits_cache,
  output [2:0] io_mmio_axi_0_aw_bits_prot,
  output [3:0] io_mmio_axi_0_aw_bits_qos,
  output [3:0] io_mmio_axi_0_aw_bits_region,
  output [4:0] io_mmio_axi_0_aw_bits_id,
  output  io_mmio_axi_0_aw_bits_user,
  input   io_mmio_axi_0_w_ready,
  output  io_mmio_axi_0_w_valid,
  output [63:0] io_mmio_axi_0_w_bits_data,
  output  io_mmio_axi_0_w_bits_last,
  output [4:0] io_mmio_axi_0_w_bits_id,
  output [7:0] io_mmio_axi_0_w_bits_strb,
  output  io_mmio_axi_0_w_bits_user,
  output  io_mmio_axi_0_b_ready,
  input   io_mmio_axi_0_b_valid,
  input  [1:0] io_mmio_axi_0_b_bits_resp,
  input  [4:0] io_mmio_axi_0_b_bits_id,
  input   io_mmio_axi_0_b_bits_user,
  input   io_mmio_axi_0_ar_ready,
  output  io_mmio_axi_0_ar_valid,
  output [31:0] io_mmio_axi_0_ar_bits_addr,
  output [7:0] io_mmio_axi_0_ar_bits_len,
  output [2:0] io_mmio_axi_0_ar_bits_size,
  output [1:0] io_mmio_axi_0_ar_bits_burst,
  output  io_mmio_axi_0_ar_bits_lock,
  output [3:0] io_mmio_axi_0_ar_bits_cache,
  output [2:0] io_mmio_axi_0_ar_bits_prot,
  output [3:0] io_mmio_axi_0_ar_bits_qos,
  output [3:0] io_mmio_axi_0_ar_bits_region,
  output [4:0] io_mmio_axi_0_ar_bits_id,
  output  io_mmio_axi_0_ar_bits_user,
  output  io_mmio_axi_0_r_ready,
  input   io_mmio_axi_0_r_valid,
  input  [1:0] io_mmio_axi_0_r_bits_resp,
  input  [63:0] io_mmio_axi_0_r_bits_data,
  input   io_mmio_axi_0_r_bits_last,
  input  [4:0] io_mmio_axi_0_r_bits_id,
  input   io_mmio_axi_0_r_bits_user,
  output  io_debug_req_ready,
  input   io_debug_req_valid,
  input  [4:0] io_debug_req_bits_addr,
  input  [1:0] io_debug_req_bits_op,
  input  [33:0] io_debug_req_bits_data,
  input   io_debug_resp_ready,
  output  io_debug_resp_valid,
  output [1:0] io_debug_resp_bits_resp,
  output [33:0] io_debug_resp_bits_data
);
//<CJ> RESET_VECTOR_ADDR
  parameter RESET_VECTOR_ADDR = 60000000;

  wire  tileResets_0;
  wire  RocketTile_1_clk;
  wire  RocketTile_1_reset;
  wire  RocketTile_1_io_cached_0_acquire_ready;
  wire  RocketTile_1_io_cached_0_acquire_valid;
  wire [25:0] RocketTile_1_io_cached_0_acquire_bits_addr_block;
  wire  RocketTile_1_io_cached_0_acquire_bits_client_xact_id;
  wire [2:0] RocketTile_1_io_cached_0_acquire_bits_addr_beat;
  wire  RocketTile_1_io_cached_0_acquire_bits_is_builtin_type;
  wire [2:0] RocketTile_1_io_cached_0_acquire_bits_a_type;
  wire [11:0] RocketTile_1_io_cached_0_acquire_bits_union;
  wire [63:0] RocketTile_1_io_cached_0_acquire_bits_data;
  wire  RocketTile_1_io_cached_0_probe_ready;
  wire  RocketTile_1_io_cached_0_probe_valid;
  wire [25:0] RocketTile_1_io_cached_0_probe_bits_addr_block;
  wire [1:0] RocketTile_1_io_cached_0_probe_bits_p_type;
  wire  RocketTile_1_io_cached_0_release_ready;
  wire  RocketTile_1_io_cached_0_release_valid;
  wire [2:0] RocketTile_1_io_cached_0_release_bits_addr_beat;
  wire [25:0] RocketTile_1_io_cached_0_release_bits_addr_block;
  wire  RocketTile_1_io_cached_0_release_bits_client_xact_id;
  wire  RocketTile_1_io_cached_0_release_bits_voluntary;
  wire [2:0] RocketTile_1_io_cached_0_release_bits_r_type;
  wire [63:0] RocketTile_1_io_cached_0_release_bits_data;
  wire  RocketTile_1_io_cached_0_grant_ready;
  wire  RocketTile_1_io_cached_0_grant_valid;
  wire [2:0] RocketTile_1_io_cached_0_grant_bits_addr_beat;
  wire  RocketTile_1_io_cached_0_grant_bits_client_xact_id;
  wire [1:0] RocketTile_1_io_cached_0_grant_bits_manager_xact_id;
  wire  RocketTile_1_io_cached_0_grant_bits_is_builtin_type;
  wire [3:0] RocketTile_1_io_cached_0_grant_bits_g_type;
  wire [63:0] RocketTile_1_io_cached_0_grant_bits_data;
  wire  RocketTile_1_io_cached_0_grant_bits_manager_id;
  wire  RocketTile_1_io_cached_0_finish_ready;
  wire  RocketTile_1_io_cached_0_finish_valid;
  wire [1:0] RocketTile_1_io_cached_0_finish_bits_manager_xact_id;
  wire  RocketTile_1_io_cached_0_finish_bits_manager_id;
  wire  RocketTile_1_io_uncached_0_acquire_ready;
  wire  RocketTile_1_io_uncached_0_acquire_valid;
  wire [25:0] RocketTile_1_io_uncached_0_acquire_bits_addr_block;
  wire  RocketTile_1_io_uncached_0_acquire_bits_client_xact_id;
  wire [2:0] RocketTile_1_io_uncached_0_acquire_bits_addr_beat;
  wire  RocketTile_1_io_uncached_0_acquire_bits_is_builtin_type;
  wire [2:0] RocketTile_1_io_uncached_0_acquire_bits_a_type;
  wire [11:0] RocketTile_1_io_uncached_0_acquire_bits_union;
  wire [63:0] RocketTile_1_io_uncached_0_acquire_bits_data;
  wire  RocketTile_1_io_uncached_0_grant_ready;
  wire  RocketTile_1_io_uncached_0_grant_valid;
  wire [2:0] RocketTile_1_io_uncached_0_grant_bits_addr_beat;
  wire  RocketTile_1_io_uncached_0_grant_bits_client_xact_id;
  wire [1:0] RocketTile_1_io_uncached_0_grant_bits_manager_xact_id;
  wire  RocketTile_1_io_uncached_0_grant_bits_is_builtin_type;
  wire [3:0] RocketTile_1_io_uncached_0_grant_bits_g_type;
  wire [63:0] RocketTile_1_io_uncached_0_grant_bits_data;
  wire  RocketTile_1_io_prci_reset;
  wire  RocketTile_1_io_prci_id;
  wire  RocketTile_1_io_prci_interrupts_meip;
  wire  RocketTile_1_io_prci_interrupts_seip;
  wire  RocketTile_1_io_prci_interrupts_debug;
  wire  RocketTile_1_io_prci_interrupts_mtip;
  wire  RocketTile_1_io_prci_interrupts_msip;
  wire  uncore_clk;
  wire  uncore_reset;
  wire  uncore_io_mem_axi_0_aw_ready;
  wire  uncore_io_mem_axi_0_aw_valid;
  wire [31:0] uncore_io_mem_axi_0_aw_bits_addr;
  wire [7:0] uncore_io_mem_axi_0_aw_bits_len;
  wire [2:0] uncore_io_mem_axi_0_aw_bits_size;
  wire [1:0] uncore_io_mem_axi_0_aw_bits_burst;
  wire  uncore_io_mem_axi_0_aw_bits_lock;
  wire [3:0] uncore_io_mem_axi_0_aw_bits_cache;
  wire [2:0] uncore_io_mem_axi_0_aw_bits_prot;
  wire [3:0] uncore_io_mem_axi_0_aw_bits_qos;
  wire [3:0] uncore_io_mem_axi_0_aw_bits_region;
  wire [4:0] uncore_io_mem_axi_0_aw_bits_id;
  wire  uncore_io_mem_axi_0_aw_bits_user;
  wire  uncore_io_mem_axi_0_w_ready;
  wire  uncore_io_mem_axi_0_w_valid;
  wire [63:0] uncore_io_mem_axi_0_w_bits_data;
  wire  uncore_io_mem_axi_0_w_bits_last;
  wire [4:0] uncore_io_mem_axi_0_w_bits_id;
  wire [7:0] uncore_io_mem_axi_0_w_bits_strb;
  wire  uncore_io_mem_axi_0_w_bits_user;
  wire  uncore_io_mem_axi_0_b_ready;
  wire  uncore_io_mem_axi_0_b_valid;
  wire [1:0] uncore_io_mem_axi_0_b_bits_resp;
  wire [4:0] uncore_io_mem_axi_0_b_bits_id;
  wire  uncore_io_mem_axi_0_b_bits_user;
  wire  uncore_io_mem_axi_0_ar_ready;
  wire  uncore_io_mem_axi_0_ar_valid;
  wire [31:0] uncore_io_mem_axi_0_ar_bits_addr;
  wire [7:0] uncore_io_mem_axi_0_ar_bits_len;
  wire [2:0] uncore_io_mem_axi_0_ar_bits_size;
  wire [1:0] uncore_io_mem_axi_0_ar_bits_burst;
  wire  uncore_io_mem_axi_0_ar_bits_lock;
  wire [3:0] uncore_io_mem_axi_0_ar_bits_cache;
  wire [2:0] uncore_io_mem_axi_0_ar_bits_prot;
  wire [3:0] uncore_io_mem_axi_0_ar_bits_qos;
  wire [3:0] uncore_io_mem_axi_0_ar_bits_region;
  wire [4:0] uncore_io_mem_axi_0_ar_bits_id;
  wire  uncore_io_mem_axi_0_ar_bits_user;
  wire  uncore_io_mem_axi_0_r_ready;
  wire  uncore_io_mem_axi_0_r_valid;
  wire [1:0] uncore_io_mem_axi_0_r_bits_resp;
  wire [63:0] uncore_io_mem_axi_0_r_bits_data;
  wire  uncore_io_mem_axi_0_r_bits_last;
  wire [4:0] uncore_io_mem_axi_0_r_bits_id;
  wire  uncore_io_mem_axi_0_r_bits_user;
  wire  uncore_io_tiles_cached_0_acquire_ready;
  wire  uncore_io_tiles_cached_0_acquire_valid;
  wire [25:0] uncore_io_tiles_cached_0_acquire_bits_addr_block;
  wire  uncore_io_tiles_cached_0_acquire_bits_client_xact_id;
  wire [2:0] uncore_io_tiles_cached_0_acquire_bits_addr_beat;
  wire  uncore_io_tiles_cached_0_acquire_bits_is_builtin_type;
  wire [2:0] uncore_io_tiles_cached_0_acquire_bits_a_type;
  wire [11:0] uncore_io_tiles_cached_0_acquire_bits_union;
  wire [63:0] uncore_io_tiles_cached_0_acquire_bits_data;
  wire  uncore_io_tiles_cached_0_probe_ready;
  wire  uncore_io_tiles_cached_0_probe_valid;
  wire [25:0] uncore_io_tiles_cached_0_probe_bits_addr_block;
  wire [1:0] uncore_io_tiles_cached_0_probe_bits_p_type;
  wire  uncore_io_tiles_cached_0_release_ready;
  wire  uncore_io_tiles_cached_0_release_valid;
  wire [2:0] uncore_io_tiles_cached_0_release_bits_addr_beat;
  wire [25:0] uncore_io_tiles_cached_0_release_bits_addr_block;
  wire  uncore_io_tiles_cached_0_release_bits_client_xact_id;
  wire  uncore_io_tiles_cached_0_release_bits_voluntary;
  wire [2:0] uncore_io_tiles_cached_0_release_bits_r_type;
  wire [63:0] uncore_io_tiles_cached_0_release_bits_data;
  wire  uncore_io_tiles_cached_0_grant_ready;
  wire  uncore_io_tiles_cached_0_grant_valid;
  wire [2:0] uncore_io_tiles_cached_0_grant_bits_addr_beat;
  wire  uncore_io_tiles_cached_0_grant_bits_client_xact_id;
  wire [1:0] uncore_io_tiles_cached_0_grant_bits_manager_xact_id;
  wire  uncore_io_tiles_cached_0_grant_bits_is_builtin_type;
  wire [3:0] uncore_io_tiles_cached_0_grant_bits_g_type;
  wire [63:0] uncore_io_tiles_cached_0_grant_bits_data;
  wire  uncore_io_tiles_cached_0_grant_bits_manager_id;
  wire  uncore_io_tiles_cached_0_finish_ready;
  wire  uncore_io_tiles_cached_0_finish_valid;
  wire [1:0] uncore_io_tiles_cached_0_finish_bits_manager_xact_id;
  wire  uncore_io_tiles_cached_0_finish_bits_manager_id;
  wire  uncore_io_tiles_uncached_0_acquire_ready;
  wire  uncore_io_tiles_uncached_0_acquire_valid;
  wire [25:0] uncore_io_tiles_uncached_0_acquire_bits_addr_block;
  wire  uncore_io_tiles_uncached_0_acquire_bits_client_xact_id;
  wire [2:0] uncore_io_tiles_uncached_0_acquire_bits_addr_beat;
  wire  uncore_io_tiles_uncached_0_acquire_bits_is_builtin_type;
  wire [2:0] uncore_io_tiles_uncached_0_acquire_bits_a_type;
  wire [11:0] uncore_io_tiles_uncached_0_acquire_bits_union;
  wire [63:0] uncore_io_tiles_uncached_0_acquire_bits_data;
  wire  uncore_io_tiles_uncached_0_grant_ready;
  wire  uncore_io_tiles_uncached_0_grant_valid;
  wire [2:0] uncore_io_tiles_uncached_0_grant_bits_addr_beat;
  wire  uncore_io_tiles_uncached_0_grant_bits_client_xact_id;
  wire [1:0] uncore_io_tiles_uncached_0_grant_bits_manager_xact_id;
  wire  uncore_io_tiles_uncached_0_grant_bits_is_builtin_type;
  wire [3:0] uncore_io_tiles_uncached_0_grant_bits_g_type;
  wire [63:0] uncore_io_tiles_uncached_0_grant_bits_data;
  wire  uncore_io_prci_0_reset;
  wire  uncore_io_prci_0_id;
  wire  uncore_io_prci_0_interrupts_meip;
  wire  uncore_io_prci_0_interrupts_seip;
  wire  uncore_io_prci_0_interrupts_debug;
  wire  uncore_io_prci_0_interrupts_mtip;
  wire  uncore_io_prci_0_interrupts_msip;
  wire  uncore_io_mmio_axi_0_aw_ready;
  wire  uncore_io_mmio_axi_0_aw_valid;
  wire [31:0] uncore_io_mmio_axi_0_aw_bits_addr;
  wire [7:0] uncore_io_mmio_axi_0_aw_bits_len;
  wire [2:0] uncore_io_mmio_axi_0_aw_bits_size;
  wire [1:0] uncore_io_mmio_axi_0_aw_bits_burst;
  wire  uncore_io_mmio_axi_0_aw_bits_lock;
  wire [3:0] uncore_io_mmio_axi_0_aw_bits_cache;
  wire [2:0] uncore_io_mmio_axi_0_aw_bits_prot;
  wire [3:0] uncore_io_mmio_axi_0_aw_bits_qos;
  wire [3:0] uncore_io_mmio_axi_0_aw_bits_region;
  wire [4:0] uncore_io_mmio_axi_0_aw_bits_id;
  wire  uncore_io_mmio_axi_0_aw_bits_user;
  wire  uncore_io_mmio_axi_0_w_ready;
  wire  uncore_io_mmio_axi_0_w_valid;
  wire [63:0] uncore_io_mmio_axi_0_w_bits_data;
  wire  uncore_io_mmio_axi_0_w_bits_last;
  wire [4:0] uncore_io_mmio_axi_0_w_bits_id;
  wire [7:0] uncore_io_mmio_axi_0_w_bits_strb;
  wire  uncore_io_mmio_axi_0_w_bits_user;
  wire  uncore_io_mmio_axi_0_b_ready;
  wire  uncore_io_mmio_axi_0_b_valid;
  wire [1:0] uncore_io_mmio_axi_0_b_bits_resp;
  wire [4:0] uncore_io_mmio_axi_0_b_bits_id;
  wire  uncore_io_mmio_axi_0_b_bits_user;
  wire  uncore_io_mmio_axi_0_ar_ready;
  wire  uncore_io_mmio_axi_0_ar_valid;
  wire [31:0] uncore_io_mmio_axi_0_ar_bits_addr;
  wire [7:0] uncore_io_mmio_axi_0_ar_bits_len;
  wire [2:0] uncore_io_mmio_axi_0_ar_bits_size;
  wire [1:0] uncore_io_mmio_axi_0_ar_bits_burst;
  wire  uncore_io_mmio_axi_0_ar_bits_lock;
  wire [3:0] uncore_io_mmio_axi_0_ar_bits_cache;
  wire [2:0] uncore_io_mmio_axi_0_ar_bits_prot;
  wire [3:0] uncore_io_mmio_axi_0_ar_bits_qos;
  wire [3:0] uncore_io_mmio_axi_0_ar_bits_region;
  wire [4:0] uncore_io_mmio_axi_0_ar_bits_id;
  wire  uncore_io_mmio_axi_0_ar_bits_user;
  wire  uncore_io_mmio_axi_0_r_ready;
  wire  uncore_io_mmio_axi_0_r_valid;
  wire [1:0] uncore_io_mmio_axi_0_r_bits_resp;
  wire [63:0] uncore_io_mmio_axi_0_r_bits_data;
  wire  uncore_io_mmio_axi_0_r_bits_last;
  wire [4:0] uncore_io_mmio_axi_0_r_bits_id;
  wire  uncore_io_mmio_axi_0_r_bits_user;
  wire  uncore_io_interrupts_0;
  wire  uncore_io_interrupts_1;
  wire  uncore_io_interrupts_2;
  wire  uncore_io_interrupts_3;
  wire  uncore_io_interrupts_4;
  wire  uncore_io_interrupts_5;
  wire  uncore_io_interrupts_6;
  wire  uncore_io_interrupts_7;
  wire  uncore_io_interrupts_8;
  wire  uncore_io_interrupts_9;
  wire  uncore_io_interrupts_10;
  wire  uncore_io_interrupts_11;
  wire  uncore_io_interrupts_12;
  wire  uncore_io_interrupts_13;
  wire  uncore_io_interrupts_14;
  wire  uncore_io_interrupts_15;
  wire  uncore_io_interrupts_16;
  wire  uncore_io_interrupts_17;
  wire  uncore_io_interrupts_18;
  wire  uncore_io_interrupts_19;
  wire  uncore_io_interrupts_20;
  wire  uncore_io_interrupts_21;
  wire  uncore_io_interrupts_22;
  wire  uncore_io_interrupts_23;
  wire  uncore_io_interrupts_24;
  wire  uncore_io_interrupts_25;
  wire  uncore_io_interrupts_26;
  wire  uncore_io_interrupts_27;
  wire  uncore_io_interrupts_28;
  wire  uncore_io_interrupts_29;
  wire  uncore_io_interrupts_30;
  wire  uncore_io_debugBus_req_ready;
  wire  uncore_io_debugBus_req_valid;
  wire [4:0] uncore_io_debugBus_req_bits_addr;
  wire [1:0] uncore_io_debugBus_req_bits_op;
  wire [33:0] uncore_io_debugBus_req_bits_data;
  wire  uncore_io_debugBus_resp_ready;
  wire  uncore_io_debugBus_resp_valid;
  wire [1:0] uncore_io_debugBus_resp_bits_resp;
  wire [33:0] uncore_io_debugBus_resp_bits_data;
  
  //<CJ> RESET_VECTOR_ADDR
   defparam RocketTile_1.RESET_VECTOR_ADDR = RESET_VECTOR_ADDR;

  RocketTile RocketTile_1 (
    .clk(RocketTile_1_clk),
    .reset(RocketTile_1_reset),
    .io_cached_0_acquire_ready(RocketTile_1_io_cached_0_acquire_ready),
    .io_cached_0_acquire_valid(RocketTile_1_io_cached_0_acquire_valid),
    .io_cached_0_acquire_bits_addr_block(RocketTile_1_io_cached_0_acquire_bits_addr_block),
    .io_cached_0_acquire_bits_client_xact_id(RocketTile_1_io_cached_0_acquire_bits_client_xact_id),
    .io_cached_0_acquire_bits_addr_beat(RocketTile_1_io_cached_0_acquire_bits_addr_beat),
    .io_cached_0_acquire_bits_is_builtin_type(RocketTile_1_io_cached_0_acquire_bits_is_builtin_type),
    .io_cached_0_acquire_bits_a_type(RocketTile_1_io_cached_0_acquire_bits_a_type),
    .io_cached_0_acquire_bits_union(RocketTile_1_io_cached_0_acquire_bits_union),
    .io_cached_0_acquire_bits_data(RocketTile_1_io_cached_0_acquire_bits_data),
    .io_cached_0_probe_ready(RocketTile_1_io_cached_0_probe_ready),
    .io_cached_0_probe_valid(RocketTile_1_io_cached_0_probe_valid),
    .io_cached_0_probe_bits_addr_block(RocketTile_1_io_cached_0_probe_bits_addr_block),
    .io_cached_0_probe_bits_p_type(RocketTile_1_io_cached_0_probe_bits_p_type),
    .io_cached_0_release_ready(RocketTile_1_io_cached_0_release_ready),
    .io_cached_0_release_valid(RocketTile_1_io_cached_0_release_valid),
    .io_cached_0_release_bits_addr_beat(RocketTile_1_io_cached_0_release_bits_addr_beat),
    .io_cached_0_release_bits_addr_block(RocketTile_1_io_cached_0_release_bits_addr_block),
    .io_cached_0_release_bits_client_xact_id(RocketTile_1_io_cached_0_release_bits_client_xact_id),
    .io_cached_0_release_bits_voluntary(RocketTile_1_io_cached_0_release_bits_voluntary),
    .io_cached_0_release_bits_r_type(RocketTile_1_io_cached_0_release_bits_r_type),
    .io_cached_0_release_bits_data(RocketTile_1_io_cached_0_release_bits_data),
    .io_cached_0_grant_ready(RocketTile_1_io_cached_0_grant_ready),
    .io_cached_0_grant_valid(RocketTile_1_io_cached_0_grant_valid),
    .io_cached_0_grant_bits_addr_beat(RocketTile_1_io_cached_0_grant_bits_addr_beat),
    .io_cached_0_grant_bits_client_xact_id(RocketTile_1_io_cached_0_grant_bits_client_xact_id),
    .io_cached_0_grant_bits_manager_xact_id(RocketTile_1_io_cached_0_grant_bits_manager_xact_id),
    .io_cached_0_grant_bits_is_builtin_type(RocketTile_1_io_cached_0_grant_bits_is_builtin_type),
    .io_cached_0_grant_bits_g_type(RocketTile_1_io_cached_0_grant_bits_g_type),
    .io_cached_0_grant_bits_data(RocketTile_1_io_cached_0_grant_bits_data),
    .io_cached_0_grant_bits_manager_id(RocketTile_1_io_cached_0_grant_bits_manager_id),
    .io_cached_0_finish_ready(RocketTile_1_io_cached_0_finish_ready),
    .io_cached_0_finish_valid(RocketTile_1_io_cached_0_finish_valid),
    .io_cached_0_finish_bits_manager_xact_id(RocketTile_1_io_cached_0_finish_bits_manager_xact_id),
    .io_cached_0_finish_bits_manager_id(RocketTile_1_io_cached_0_finish_bits_manager_id),
    .io_uncached_0_acquire_ready(RocketTile_1_io_uncached_0_acquire_ready),
    .io_uncached_0_acquire_valid(RocketTile_1_io_uncached_0_acquire_valid),
    .io_uncached_0_acquire_bits_addr_block(RocketTile_1_io_uncached_0_acquire_bits_addr_block),
    .io_uncached_0_acquire_bits_client_xact_id(RocketTile_1_io_uncached_0_acquire_bits_client_xact_id),
    .io_uncached_0_acquire_bits_addr_beat(RocketTile_1_io_uncached_0_acquire_bits_addr_beat),
    .io_uncached_0_acquire_bits_is_builtin_type(RocketTile_1_io_uncached_0_acquire_bits_is_builtin_type),
    .io_uncached_0_acquire_bits_a_type(RocketTile_1_io_uncached_0_acquire_bits_a_type),
    .io_uncached_0_acquire_bits_union(RocketTile_1_io_uncached_0_acquire_bits_union),
    .io_uncached_0_acquire_bits_data(RocketTile_1_io_uncached_0_acquire_bits_data),
    .io_uncached_0_grant_ready(RocketTile_1_io_uncached_0_grant_ready),
    .io_uncached_0_grant_valid(RocketTile_1_io_uncached_0_grant_valid),
    .io_uncached_0_grant_bits_addr_beat(RocketTile_1_io_uncached_0_grant_bits_addr_beat),
    .io_uncached_0_grant_bits_client_xact_id(RocketTile_1_io_uncached_0_grant_bits_client_xact_id),
    .io_uncached_0_grant_bits_manager_xact_id(RocketTile_1_io_uncached_0_grant_bits_manager_xact_id),
    .io_uncached_0_grant_bits_is_builtin_type(RocketTile_1_io_uncached_0_grant_bits_is_builtin_type),
    .io_uncached_0_grant_bits_g_type(RocketTile_1_io_uncached_0_grant_bits_g_type),
    .io_uncached_0_grant_bits_data(RocketTile_1_io_uncached_0_grant_bits_data),
    .io_prci_reset(RocketTile_1_io_prci_reset),
    .io_prci_id(RocketTile_1_io_prci_id),
    .io_prci_interrupts_meip(RocketTile_1_io_prci_interrupts_meip),
    .io_prci_interrupts_seip(RocketTile_1_io_prci_interrupts_seip),
    .io_prci_interrupts_debug(RocketTile_1_io_prci_interrupts_debug),
    .io_prci_interrupts_mtip(RocketTile_1_io_prci_interrupts_mtip),
    .io_prci_interrupts_msip(RocketTile_1_io_prci_interrupts_msip)
  );
  Uncore uncore (
    .clk(uncore_clk),
    .reset(uncore_reset),
    .io_mem_axi_0_aw_ready(uncore_io_mem_axi_0_aw_ready),
    .io_mem_axi_0_aw_valid(uncore_io_mem_axi_0_aw_valid),
    .io_mem_axi_0_aw_bits_addr(uncore_io_mem_axi_0_aw_bits_addr),
    .io_mem_axi_0_aw_bits_len(uncore_io_mem_axi_0_aw_bits_len),
    .io_mem_axi_0_aw_bits_size(uncore_io_mem_axi_0_aw_bits_size),
    .io_mem_axi_0_aw_bits_burst(uncore_io_mem_axi_0_aw_bits_burst),
    .io_mem_axi_0_aw_bits_lock(uncore_io_mem_axi_0_aw_bits_lock),
    .io_mem_axi_0_aw_bits_cache(uncore_io_mem_axi_0_aw_bits_cache),
    .io_mem_axi_0_aw_bits_prot(uncore_io_mem_axi_0_aw_bits_prot),
    .io_mem_axi_0_aw_bits_qos(uncore_io_mem_axi_0_aw_bits_qos),
    .io_mem_axi_0_aw_bits_region(uncore_io_mem_axi_0_aw_bits_region),
    .io_mem_axi_0_aw_bits_id(uncore_io_mem_axi_0_aw_bits_id),
    .io_mem_axi_0_aw_bits_user(uncore_io_mem_axi_0_aw_bits_user),
    .io_mem_axi_0_w_ready(uncore_io_mem_axi_0_w_ready),
    .io_mem_axi_0_w_valid(uncore_io_mem_axi_0_w_valid),
    .io_mem_axi_0_w_bits_data(uncore_io_mem_axi_0_w_bits_data),
    .io_mem_axi_0_w_bits_last(uncore_io_mem_axi_0_w_bits_last),
    .io_mem_axi_0_w_bits_id(uncore_io_mem_axi_0_w_bits_id),
    .io_mem_axi_0_w_bits_strb(uncore_io_mem_axi_0_w_bits_strb),
    .io_mem_axi_0_w_bits_user(uncore_io_mem_axi_0_w_bits_user),
    .io_mem_axi_0_b_ready(uncore_io_mem_axi_0_b_ready),
    .io_mem_axi_0_b_valid(uncore_io_mem_axi_0_b_valid),
    .io_mem_axi_0_b_bits_resp(uncore_io_mem_axi_0_b_bits_resp),
    .io_mem_axi_0_b_bits_id(uncore_io_mem_axi_0_b_bits_id),
    .io_mem_axi_0_b_bits_user(uncore_io_mem_axi_0_b_bits_user),
    .io_mem_axi_0_ar_ready(uncore_io_mem_axi_0_ar_ready),
    .io_mem_axi_0_ar_valid(uncore_io_mem_axi_0_ar_valid),
    .io_mem_axi_0_ar_bits_addr(uncore_io_mem_axi_0_ar_bits_addr),
    .io_mem_axi_0_ar_bits_len(uncore_io_mem_axi_0_ar_bits_len),
    .io_mem_axi_0_ar_bits_size(uncore_io_mem_axi_0_ar_bits_size),
    .io_mem_axi_0_ar_bits_burst(uncore_io_mem_axi_0_ar_bits_burst),
    .io_mem_axi_0_ar_bits_lock(uncore_io_mem_axi_0_ar_bits_lock),
    .io_mem_axi_0_ar_bits_cache(uncore_io_mem_axi_0_ar_bits_cache),
    .io_mem_axi_0_ar_bits_prot(uncore_io_mem_axi_0_ar_bits_prot),
    .io_mem_axi_0_ar_bits_qos(uncore_io_mem_axi_0_ar_bits_qos),
    .io_mem_axi_0_ar_bits_region(uncore_io_mem_axi_0_ar_bits_region),
    .io_mem_axi_0_ar_bits_id(uncore_io_mem_axi_0_ar_bits_id),
    .io_mem_axi_0_ar_bits_user(uncore_io_mem_axi_0_ar_bits_user),
    .io_mem_axi_0_r_ready(uncore_io_mem_axi_0_r_ready),
    .io_mem_axi_0_r_valid(uncore_io_mem_axi_0_r_valid),
    .io_mem_axi_0_r_bits_resp(uncore_io_mem_axi_0_r_bits_resp),
    .io_mem_axi_0_r_bits_data(uncore_io_mem_axi_0_r_bits_data),
    .io_mem_axi_0_r_bits_last(uncore_io_mem_axi_0_r_bits_last),
    .io_mem_axi_0_r_bits_id(uncore_io_mem_axi_0_r_bits_id),
    .io_mem_axi_0_r_bits_user(uncore_io_mem_axi_0_r_bits_user),
    .io_tiles_cached_0_acquire_ready(uncore_io_tiles_cached_0_acquire_ready),
    .io_tiles_cached_0_acquire_valid(uncore_io_tiles_cached_0_acquire_valid),
    .io_tiles_cached_0_acquire_bits_addr_block(uncore_io_tiles_cached_0_acquire_bits_addr_block),
    .io_tiles_cached_0_acquire_bits_client_xact_id(uncore_io_tiles_cached_0_acquire_bits_client_xact_id),
    .io_tiles_cached_0_acquire_bits_addr_beat(uncore_io_tiles_cached_0_acquire_bits_addr_beat),
    .io_tiles_cached_0_acquire_bits_is_builtin_type(uncore_io_tiles_cached_0_acquire_bits_is_builtin_type),
    .io_tiles_cached_0_acquire_bits_a_type(uncore_io_tiles_cached_0_acquire_bits_a_type),
    .io_tiles_cached_0_acquire_bits_union(uncore_io_tiles_cached_0_acquire_bits_union),
    .io_tiles_cached_0_acquire_bits_data(uncore_io_tiles_cached_0_acquire_bits_data),
    .io_tiles_cached_0_probe_ready(uncore_io_tiles_cached_0_probe_ready),
    .io_tiles_cached_0_probe_valid(uncore_io_tiles_cached_0_probe_valid),
    .io_tiles_cached_0_probe_bits_addr_block(uncore_io_tiles_cached_0_probe_bits_addr_block),
    .io_tiles_cached_0_probe_bits_p_type(uncore_io_tiles_cached_0_probe_bits_p_type),
    .io_tiles_cached_0_release_ready(uncore_io_tiles_cached_0_release_ready),
    .io_tiles_cached_0_release_valid(uncore_io_tiles_cached_0_release_valid),
    .io_tiles_cached_0_release_bits_addr_beat(uncore_io_tiles_cached_0_release_bits_addr_beat),
    .io_tiles_cached_0_release_bits_addr_block(uncore_io_tiles_cached_0_release_bits_addr_block),
    .io_tiles_cached_0_release_bits_client_xact_id(uncore_io_tiles_cached_0_release_bits_client_xact_id),
    .io_tiles_cached_0_release_bits_voluntary(uncore_io_tiles_cached_0_release_bits_voluntary),
    .io_tiles_cached_0_release_bits_r_type(uncore_io_tiles_cached_0_release_bits_r_type),
    .io_tiles_cached_0_release_bits_data(uncore_io_tiles_cached_0_release_bits_data),
    .io_tiles_cached_0_grant_ready(uncore_io_tiles_cached_0_grant_ready),
    .io_tiles_cached_0_grant_valid(uncore_io_tiles_cached_0_grant_valid),
    .io_tiles_cached_0_grant_bits_addr_beat(uncore_io_tiles_cached_0_grant_bits_addr_beat),
    .io_tiles_cached_0_grant_bits_client_xact_id(uncore_io_tiles_cached_0_grant_bits_client_xact_id),
    .io_tiles_cached_0_grant_bits_manager_xact_id(uncore_io_tiles_cached_0_grant_bits_manager_xact_id),
    .io_tiles_cached_0_grant_bits_is_builtin_type(uncore_io_tiles_cached_0_grant_bits_is_builtin_type),
    .io_tiles_cached_0_grant_bits_g_type(uncore_io_tiles_cached_0_grant_bits_g_type),
    .io_tiles_cached_0_grant_bits_data(uncore_io_tiles_cached_0_grant_bits_data),
    .io_tiles_cached_0_grant_bits_manager_id(uncore_io_tiles_cached_0_grant_bits_manager_id),
    .io_tiles_cached_0_finish_ready(uncore_io_tiles_cached_0_finish_ready),
    .io_tiles_cached_0_finish_valid(uncore_io_tiles_cached_0_finish_valid),
    .io_tiles_cached_0_finish_bits_manager_xact_id(uncore_io_tiles_cached_0_finish_bits_manager_xact_id),
    .io_tiles_cached_0_finish_bits_manager_id(uncore_io_tiles_cached_0_finish_bits_manager_id),
    .io_tiles_uncached_0_acquire_ready(uncore_io_tiles_uncached_0_acquire_ready),
    .io_tiles_uncached_0_acquire_valid(uncore_io_tiles_uncached_0_acquire_valid),
    .io_tiles_uncached_0_acquire_bits_addr_block(uncore_io_tiles_uncached_0_acquire_bits_addr_block),
    .io_tiles_uncached_0_acquire_bits_client_xact_id(uncore_io_tiles_uncached_0_acquire_bits_client_xact_id),
    .io_tiles_uncached_0_acquire_bits_addr_beat(uncore_io_tiles_uncached_0_acquire_bits_addr_beat),
    .io_tiles_uncached_0_acquire_bits_is_builtin_type(uncore_io_tiles_uncached_0_acquire_bits_is_builtin_type),
    .io_tiles_uncached_0_acquire_bits_a_type(uncore_io_tiles_uncached_0_acquire_bits_a_type),
    .io_tiles_uncached_0_acquire_bits_union(uncore_io_tiles_uncached_0_acquire_bits_union),
    .io_tiles_uncached_0_acquire_bits_data(uncore_io_tiles_uncached_0_acquire_bits_data),
    .io_tiles_uncached_0_grant_ready(uncore_io_tiles_uncached_0_grant_ready),
    .io_tiles_uncached_0_grant_valid(uncore_io_tiles_uncached_0_grant_valid),
    .io_tiles_uncached_0_grant_bits_addr_beat(uncore_io_tiles_uncached_0_grant_bits_addr_beat),
    .io_tiles_uncached_0_grant_bits_client_xact_id(uncore_io_tiles_uncached_0_grant_bits_client_xact_id),
    .io_tiles_uncached_0_grant_bits_manager_xact_id(uncore_io_tiles_uncached_0_grant_bits_manager_xact_id),
    .io_tiles_uncached_0_grant_bits_is_builtin_type(uncore_io_tiles_uncached_0_grant_bits_is_builtin_type),
    .io_tiles_uncached_0_grant_bits_g_type(uncore_io_tiles_uncached_0_grant_bits_g_type),
    .io_tiles_uncached_0_grant_bits_data(uncore_io_tiles_uncached_0_grant_bits_data),
    .io_prci_0_reset(uncore_io_prci_0_reset),
    .io_prci_0_id(uncore_io_prci_0_id),
    .io_prci_0_interrupts_meip(uncore_io_prci_0_interrupts_meip),
    .io_prci_0_interrupts_seip(uncore_io_prci_0_interrupts_seip),
    .io_prci_0_interrupts_debug(uncore_io_prci_0_interrupts_debug),
    .io_prci_0_interrupts_mtip(uncore_io_prci_0_interrupts_mtip),
    .io_prci_0_interrupts_msip(uncore_io_prci_0_interrupts_msip),
    .io_mmio_axi_0_aw_ready(uncore_io_mmio_axi_0_aw_ready),
    .io_mmio_axi_0_aw_valid(uncore_io_mmio_axi_0_aw_valid),
    .io_mmio_axi_0_aw_bits_addr(uncore_io_mmio_axi_0_aw_bits_addr),
    .io_mmio_axi_0_aw_bits_len(uncore_io_mmio_axi_0_aw_bits_len),
    .io_mmio_axi_0_aw_bits_size(uncore_io_mmio_axi_0_aw_bits_size),
    .io_mmio_axi_0_aw_bits_burst(uncore_io_mmio_axi_0_aw_bits_burst),
    .io_mmio_axi_0_aw_bits_lock(uncore_io_mmio_axi_0_aw_bits_lock),
    .io_mmio_axi_0_aw_bits_cache(uncore_io_mmio_axi_0_aw_bits_cache),
    .io_mmio_axi_0_aw_bits_prot(uncore_io_mmio_axi_0_aw_bits_prot),
    .io_mmio_axi_0_aw_bits_qos(uncore_io_mmio_axi_0_aw_bits_qos),
    .io_mmio_axi_0_aw_bits_region(uncore_io_mmio_axi_0_aw_bits_region),
    .io_mmio_axi_0_aw_bits_id(uncore_io_mmio_axi_0_aw_bits_id),
    .io_mmio_axi_0_aw_bits_user(uncore_io_mmio_axi_0_aw_bits_user),
    .io_mmio_axi_0_w_ready(uncore_io_mmio_axi_0_w_ready),
    .io_mmio_axi_0_w_valid(uncore_io_mmio_axi_0_w_valid),
    .io_mmio_axi_0_w_bits_data(uncore_io_mmio_axi_0_w_bits_data),
    .io_mmio_axi_0_w_bits_last(uncore_io_mmio_axi_0_w_bits_last),
    .io_mmio_axi_0_w_bits_id(uncore_io_mmio_axi_0_w_bits_id),
    .io_mmio_axi_0_w_bits_strb(uncore_io_mmio_axi_0_w_bits_strb),
    .io_mmio_axi_0_w_bits_user(uncore_io_mmio_axi_0_w_bits_user),
    .io_mmio_axi_0_b_ready(uncore_io_mmio_axi_0_b_ready),
    .io_mmio_axi_0_b_valid(uncore_io_mmio_axi_0_b_valid),
    .io_mmio_axi_0_b_bits_resp(uncore_io_mmio_axi_0_b_bits_resp),
    .io_mmio_axi_0_b_bits_id(uncore_io_mmio_axi_0_b_bits_id),
    .io_mmio_axi_0_b_bits_user(uncore_io_mmio_axi_0_b_bits_user),
    .io_mmio_axi_0_ar_ready(uncore_io_mmio_axi_0_ar_ready),
    .io_mmio_axi_0_ar_valid(uncore_io_mmio_axi_0_ar_valid),
    .io_mmio_axi_0_ar_bits_addr(uncore_io_mmio_axi_0_ar_bits_addr),
    .io_mmio_axi_0_ar_bits_len(uncore_io_mmio_axi_0_ar_bits_len),
    .io_mmio_axi_0_ar_bits_size(uncore_io_mmio_axi_0_ar_bits_size),
    .io_mmio_axi_0_ar_bits_burst(uncore_io_mmio_axi_0_ar_bits_burst),
    .io_mmio_axi_0_ar_bits_lock(uncore_io_mmio_axi_0_ar_bits_lock),
    .io_mmio_axi_0_ar_bits_cache(uncore_io_mmio_axi_0_ar_bits_cache),
    .io_mmio_axi_0_ar_bits_prot(uncore_io_mmio_axi_0_ar_bits_prot),
    .io_mmio_axi_0_ar_bits_qos(uncore_io_mmio_axi_0_ar_bits_qos),
    .io_mmio_axi_0_ar_bits_region(uncore_io_mmio_axi_0_ar_bits_region),
    .io_mmio_axi_0_ar_bits_id(uncore_io_mmio_axi_0_ar_bits_id),
    .io_mmio_axi_0_ar_bits_user(uncore_io_mmio_axi_0_ar_bits_user),
    .io_mmio_axi_0_r_ready(uncore_io_mmio_axi_0_r_ready),
    .io_mmio_axi_0_r_valid(uncore_io_mmio_axi_0_r_valid),
    .io_mmio_axi_0_r_bits_resp(uncore_io_mmio_axi_0_r_bits_resp),
    .io_mmio_axi_0_r_bits_data(uncore_io_mmio_axi_0_r_bits_data),
    .io_mmio_axi_0_r_bits_last(uncore_io_mmio_axi_0_r_bits_last),
    .io_mmio_axi_0_r_bits_id(uncore_io_mmio_axi_0_r_bits_id),
    .io_mmio_axi_0_r_bits_user(uncore_io_mmio_axi_0_r_bits_user),
    .io_interrupts_0(uncore_io_interrupts_0),
    .io_interrupts_1(uncore_io_interrupts_1),
    .io_interrupts_2(uncore_io_interrupts_2),
    .io_interrupts_3(uncore_io_interrupts_3),
    .io_interrupts_4(uncore_io_interrupts_4),
    .io_interrupts_5(uncore_io_interrupts_5),
    .io_interrupts_6(uncore_io_interrupts_6),
    .io_interrupts_7(uncore_io_interrupts_7),
    .io_interrupts_8(uncore_io_interrupts_8),
    .io_interrupts_9(uncore_io_interrupts_9),
    .io_interrupts_10(uncore_io_interrupts_10),
    .io_interrupts_11(uncore_io_interrupts_11),
    .io_interrupts_12(uncore_io_interrupts_12),
    .io_interrupts_13(uncore_io_interrupts_13),
    .io_interrupts_14(uncore_io_interrupts_14),
    .io_interrupts_15(uncore_io_interrupts_15),
    .io_interrupts_16(uncore_io_interrupts_16),
    .io_interrupts_17(uncore_io_interrupts_17),
    .io_interrupts_18(uncore_io_interrupts_18),
    .io_interrupts_19(uncore_io_interrupts_19),
    .io_interrupts_20(uncore_io_interrupts_20),
    .io_interrupts_21(uncore_io_interrupts_21),
    .io_interrupts_22(uncore_io_interrupts_22),
    .io_interrupts_23(uncore_io_interrupts_23),
    .io_interrupts_24(uncore_io_interrupts_24),
    .io_interrupts_25(uncore_io_interrupts_25),
    .io_interrupts_26(uncore_io_interrupts_26),
    .io_interrupts_27(uncore_io_interrupts_27),
    .io_interrupts_28(uncore_io_interrupts_28),
    .io_interrupts_29(uncore_io_interrupts_29),
    .io_interrupts_30(uncore_io_interrupts_30),
    .io_debugBus_req_ready(uncore_io_debugBus_req_ready),
    .io_debugBus_req_valid(uncore_io_debugBus_req_valid),
    .io_debugBus_req_bits_addr(uncore_io_debugBus_req_bits_addr),
    .io_debugBus_req_bits_op(uncore_io_debugBus_req_bits_op),
    .io_debugBus_req_bits_data(uncore_io_debugBus_req_bits_data),
    .io_debugBus_resp_ready(uncore_io_debugBus_resp_ready),
    .io_debugBus_resp_valid(uncore_io_debugBus_resp_valid),
    .io_debugBus_resp_bits_resp(uncore_io_debugBus_resp_bits_resp),
    .io_debugBus_resp_bits_data(uncore_io_debugBus_resp_bits_data)
  );
  assign io_mem_axi_0_aw_valid = uncore_io_mem_axi_0_aw_valid;
  assign io_mem_axi_0_aw_bits_addr = uncore_io_mem_axi_0_aw_bits_addr;
  assign io_mem_axi_0_aw_bits_len = uncore_io_mem_axi_0_aw_bits_len;
  assign io_mem_axi_0_aw_bits_size = uncore_io_mem_axi_0_aw_bits_size;
  assign io_mem_axi_0_aw_bits_burst = uncore_io_mem_axi_0_aw_bits_burst;
  assign io_mem_axi_0_aw_bits_lock = uncore_io_mem_axi_0_aw_bits_lock;
  assign io_mem_axi_0_aw_bits_cache = uncore_io_mem_axi_0_aw_bits_cache;
  assign io_mem_axi_0_aw_bits_prot = uncore_io_mem_axi_0_aw_bits_prot;
  assign io_mem_axi_0_aw_bits_qos = uncore_io_mem_axi_0_aw_bits_qos;
  assign io_mem_axi_0_aw_bits_region = uncore_io_mem_axi_0_aw_bits_region;
  assign io_mem_axi_0_aw_bits_id = uncore_io_mem_axi_0_aw_bits_id;
  assign io_mem_axi_0_aw_bits_user = uncore_io_mem_axi_0_aw_bits_user;
  assign io_mem_axi_0_w_valid = uncore_io_mem_axi_0_w_valid;
  assign io_mem_axi_0_w_bits_data = uncore_io_mem_axi_0_w_bits_data;
  assign io_mem_axi_0_w_bits_last = uncore_io_mem_axi_0_w_bits_last;
  assign io_mem_axi_0_w_bits_id = uncore_io_mem_axi_0_w_bits_id;
  assign io_mem_axi_0_w_bits_strb = uncore_io_mem_axi_0_w_bits_strb;
  assign io_mem_axi_0_w_bits_user = uncore_io_mem_axi_0_w_bits_user;
  assign io_mem_axi_0_b_ready = uncore_io_mem_axi_0_b_ready;
  assign io_mem_axi_0_ar_valid = uncore_io_mem_axi_0_ar_valid;
  assign io_mem_axi_0_ar_bits_addr = uncore_io_mem_axi_0_ar_bits_addr;
  assign io_mem_axi_0_ar_bits_len = uncore_io_mem_axi_0_ar_bits_len;
  assign io_mem_axi_0_ar_bits_size = uncore_io_mem_axi_0_ar_bits_size;
  assign io_mem_axi_0_ar_bits_burst = uncore_io_mem_axi_0_ar_bits_burst;
  assign io_mem_axi_0_ar_bits_lock = uncore_io_mem_axi_0_ar_bits_lock;
  assign io_mem_axi_0_ar_bits_cache = uncore_io_mem_axi_0_ar_bits_cache;
  assign io_mem_axi_0_ar_bits_prot = uncore_io_mem_axi_0_ar_bits_prot;
  assign io_mem_axi_0_ar_bits_qos = uncore_io_mem_axi_0_ar_bits_qos;
  assign io_mem_axi_0_ar_bits_region = uncore_io_mem_axi_0_ar_bits_region;
  assign io_mem_axi_0_ar_bits_id = uncore_io_mem_axi_0_ar_bits_id;
  assign io_mem_axi_0_ar_bits_user = uncore_io_mem_axi_0_ar_bits_user;
  assign io_mem_axi_0_r_ready = uncore_io_mem_axi_0_r_ready;
  assign io_mmio_axi_0_aw_valid = uncore_io_mmio_axi_0_aw_valid;
  assign io_mmio_axi_0_aw_bits_addr = uncore_io_mmio_axi_0_aw_bits_addr;
  assign io_mmio_axi_0_aw_bits_len = uncore_io_mmio_axi_0_aw_bits_len;
  assign io_mmio_axi_0_aw_bits_size = uncore_io_mmio_axi_0_aw_bits_size;
  assign io_mmio_axi_0_aw_bits_burst = uncore_io_mmio_axi_0_aw_bits_burst;
  assign io_mmio_axi_0_aw_bits_lock = uncore_io_mmio_axi_0_aw_bits_lock;
  assign io_mmio_axi_0_aw_bits_cache = uncore_io_mmio_axi_0_aw_bits_cache;
  assign io_mmio_axi_0_aw_bits_prot = uncore_io_mmio_axi_0_aw_bits_prot;
  assign io_mmio_axi_0_aw_bits_qos = uncore_io_mmio_axi_0_aw_bits_qos;
  assign io_mmio_axi_0_aw_bits_region = uncore_io_mmio_axi_0_aw_bits_region;
  assign io_mmio_axi_0_aw_bits_id = uncore_io_mmio_axi_0_aw_bits_id;
  assign io_mmio_axi_0_aw_bits_user = uncore_io_mmio_axi_0_aw_bits_user;
  assign io_mmio_axi_0_w_valid = uncore_io_mmio_axi_0_w_valid;
  assign io_mmio_axi_0_w_bits_data = uncore_io_mmio_axi_0_w_bits_data;
  assign io_mmio_axi_0_w_bits_last = uncore_io_mmio_axi_0_w_bits_last;
  assign io_mmio_axi_0_w_bits_id = uncore_io_mmio_axi_0_w_bits_id;
  assign io_mmio_axi_0_w_bits_strb = uncore_io_mmio_axi_0_w_bits_strb;
  assign io_mmio_axi_0_w_bits_user = uncore_io_mmio_axi_0_w_bits_user;
  assign io_mmio_axi_0_b_ready = uncore_io_mmio_axi_0_b_ready;
  assign io_mmio_axi_0_ar_valid = uncore_io_mmio_axi_0_ar_valid;
  assign io_mmio_axi_0_ar_bits_addr = uncore_io_mmio_axi_0_ar_bits_addr;
  assign io_mmio_axi_0_ar_bits_len = uncore_io_mmio_axi_0_ar_bits_len;
  assign io_mmio_axi_0_ar_bits_size = uncore_io_mmio_axi_0_ar_bits_size;
  assign io_mmio_axi_0_ar_bits_burst = uncore_io_mmio_axi_0_ar_bits_burst;
  assign io_mmio_axi_0_ar_bits_lock = uncore_io_mmio_axi_0_ar_bits_lock;
  assign io_mmio_axi_0_ar_bits_cache = uncore_io_mmio_axi_0_ar_bits_cache;
  assign io_mmio_axi_0_ar_bits_prot = uncore_io_mmio_axi_0_ar_bits_prot;
  assign io_mmio_axi_0_ar_bits_qos = uncore_io_mmio_axi_0_ar_bits_qos;
  assign io_mmio_axi_0_ar_bits_region = uncore_io_mmio_axi_0_ar_bits_region;
  assign io_mmio_axi_0_ar_bits_id = uncore_io_mmio_axi_0_ar_bits_id;
  assign io_mmio_axi_0_ar_bits_user = uncore_io_mmio_axi_0_ar_bits_user;
  assign io_mmio_axi_0_r_ready = uncore_io_mmio_axi_0_r_ready;
  assign io_debug_req_ready = uncore_io_debugBus_req_ready;
  assign io_debug_resp_valid = uncore_io_debugBus_resp_valid;
  assign io_debug_resp_bits_resp = uncore_io_debugBus_resp_bits_resp;
  assign io_debug_resp_bits_data = uncore_io_debugBus_resp_bits_data;
  assign tileResets_0 = uncore_io_prci_0_reset;
  assign RocketTile_1_clk = clk;
  assign RocketTile_1_reset = tileResets_0;
  assign RocketTile_1_io_cached_0_acquire_ready = uncore_io_tiles_cached_0_acquire_ready;
  assign RocketTile_1_io_cached_0_probe_valid = uncore_io_tiles_cached_0_probe_valid;
  assign RocketTile_1_io_cached_0_probe_bits_addr_block = uncore_io_tiles_cached_0_probe_bits_addr_block;
  assign RocketTile_1_io_cached_0_probe_bits_p_type = uncore_io_tiles_cached_0_probe_bits_p_type;
  assign RocketTile_1_io_cached_0_release_ready = uncore_io_tiles_cached_0_release_ready;
  assign RocketTile_1_io_cached_0_grant_valid = uncore_io_tiles_cached_0_grant_valid;
  assign RocketTile_1_io_cached_0_grant_bits_addr_beat = uncore_io_tiles_cached_0_grant_bits_addr_beat;
  assign RocketTile_1_io_cached_0_grant_bits_client_xact_id = uncore_io_tiles_cached_0_grant_bits_client_xact_id;
  assign RocketTile_1_io_cached_0_grant_bits_manager_xact_id = uncore_io_tiles_cached_0_grant_bits_manager_xact_id;
  assign RocketTile_1_io_cached_0_grant_bits_is_builtin_type = uncore_io_tiles_cached_0_grant_bits_is_builtin_type;
  assign RocketTile_1_io_cached_0_grant_bits_g_type = uncore_io_tiles_cached_0_grant_bits_g_type;
  assign RocketTile_1_io_cached_0_grant_bits_data = uncore_io_tiles_cached_0_grant_bits_data;
  assign RocketTile_1_io_cached_0_grant_bits_manager_id = uncore_io_tiles_cached_0_grant_bits_manager_id;
  assign RocketTile_1_io_cached_0_finish_ready = uncore_io_tiles_cached_0_finish_ready;
  assign RocketTile_1_io_uncached_0_acquire_ready = uncore_io_tiles_uncached_0_acquire_ready;
  assign RocketTile_1_io_uncached_0_grant_valid = uncore_io_tiles_uncached_0_grant_valid;
  assign RocketTile_1_io_uncached_0_grant_bits_addr_beat = uncore_io_tiles_uncached_0_grant_bits_addr_beat;
  assign RocketTile_1_io_uncached_0_grant_bits_client_xact_id = uncore_io_tiles_uncached_0_grant_bits_client_xact_id;
  assign RocketTile_1_io_uncached_0_grant_bits_manager_xact_id = uncore_io_tiles_uncached_0_grant_bits_manager_xact_id;
  assign RocketTile_1_io_uncached_0_grant_bits_is_builtin_type = uncore_io_tiles_uncached_0_grant_bits_is_builtin_type;
  assign RocketTile_1_io_uncached_0_grant_bits_g_type = uncore_io_tiles_uncached_0_grant_bits_g_type;
  assign RocketTile_1_io_uncached_0_grant_bits_data = uncore_io_tiles_uncached_0_grant_bits_data;
  assign RocketTile_1_io_prci_reset = uncore_io_prci_0_reset;
  assign RocketTile_1_io_prci_id = uncore_io_prci_0_id;
  assign RocketTile_1_io_prci_interrupts_meip = uncore_io_prci_0_interrupts_meip;
  assign RocketTile_1_io_prci_interrupts_seip = uncore_io_prci_0_interrupts_seip;
  assign RocketTile_1_io_prci_interrupts_debug = uncore_io_prci_0_interrupts_debug;
  assign RocketTile_1_io_prci_interrupts_mtip = uncore_io_prci_0_interrupts_mtip;
  assign RocketTile_1_io_prci_interrupts_msip = uncore_io_prci_0_interrupts_msip;
  assign uncore_clk = clk;
  assign uncore_reset = reset;
  assign uncore_io_mem_axi_0_aw_ready = io_mem_axi_0_aw_ready;
  assign uncore_io_mem_axi_0_w_ready = io_mem_axi_0_w_ready;
  assign uncore_io_mem_axi_0_b_valid = io_mem_axi_0_b_valid;
  assign uncore_io_mem_axi_0_b_bits_resp = io_mem_axi_0_b_bits_resp;
  assign uncore_io_mem_axi_0_b_bits_id = io_mem_axi_0_b_bits_id;
  assign uncore_io_mem_axi_0_b_bits_user = io_mem_axi_0_b_bits_user;
  assign uncore_io_mem_axi_0_ar_ready = io_mem_axi_0_ar_ready;
  assign uncore_io_mem_axi_0_r_valid = io_mem_axi_0_r_valid;
  assign uncore_io_mem_axi_0_r_bits_resp = io_mem_axi_0_r_bits_resp;
  assign uncore_io_mem_axi_0_r_bits_data = io_mem_axi_0_r_bits_data;
  assign uncore_io_mem_axi_0_r_bits_last = io_mem_axi_0_r_bits_last;
  assign uncore_io_mem_axi_0_r_bits_id = io_mem_axi_0_r_bits_id;
  assign uncore_io_mem_axi_0_r_bits_user = io_mem_axi_0_r_bits_user;
  assign uncore_io_tiles_cached_0_acquire_valid = RocketTile_1_io_cached_0_acquire_valid;
  assign uncore_io_tiles_cached_0_acquire_bits_addr_block = RocketTile_1_io_cached_0_acquire_bits_addr_block;
  assign uncore_io_tiles_cached_0_acquire_bits_client_xact_id = RocketTile_1_io_cached_0_acquire_bits_client_xact_id;
  assign uncore_io_tiles_cached_0_acquire_bits_addr_beat = RocketTile_1_io_cached_0_acquire_bits_addr_beat;
  assign uncore_io_tiles_cached_0_acquire_bits_is_builtin_type = RocketTile_1_io_cached_0_acquire_bits_is_builtin_type;
  assign uncore_io_tiles_cached_0_acquire_bits_a_type = RocketTile_1_io_cached_0_acquire_bits_a_type;
  assign uncore_io_tiles_cached_0_acquire_bits_union = RocketTile_1_io_cached_0_acquire_bits_union;
  assign uncore_io_tiles_cached_0_acquire_bits_data = RocketTile_1_io_cached_0_acquire_bits_data;
  assign uncore_io_tiles_cached_0_probe_ready = RocketTile_1_io_cached_0_probe_ready;
  assign uncore_io_tiles_cached_0_release_valid = RocketTile_1_io_cached_0_release_valid;
  assign uncore_io_tiles_cached_0_release_bits_addr_beat = RocketTile_1_io_cached_0_release_bits_addr_beat;
  assign uncore_io_tiles_cached_0_release_bits_addr_block = RocketTile_1_io_cached_0_release_bits_addr_block;
  assign uncore_io_tiles_cached_0_release_bits_client_xact_id = RocketTile_1_io_cached_0_release_bits_client_xact_id;
  assign uncore_io_tiles_cached_0_release_bits_voluntary = RocketTile_1_io_cached_0_release_bits_voluntary;
  assign uncore_io_tiles_cached_0_release_bits_r_type = RocketTile_1_io_cached_0_release_bits_r_type;
  assign uncore_io_tiles_cached_0_release_bits_data = RocketTile_1_io_cached_0_release_bits_data;
  assign uncore_io_tiles_cached_0_grant_ready = RocketTile_1_io_cached_0_grant_ready;
  assign uncore_io_tiles_cached_0_finish_valid = RocketTile_1_io_cached_0_finish_valid;
  assign uncore_io_tiles_cached_0_finish_bits_manager_xact_id = RocketTile_1_io_cached_0_finish_bits_manager_xact_id;
  assign uncore_io_tiles_cached_0_finish_bits_manager_id = RocketTile_1_io_cached_0_finish_bits_manager_id;
  assign uncore_io_tiles_uncached_0_acquire_valid = RocketTile_1_io_uncached_0_acquire_valid;
  assign uncore_io_tiles_uncached_0_acquire_bits_addr_block = RocketTile_1_io_uncached_0_acquire_bits_addr_block;
  assign uncore_io_tiles_uncached_0_acquire_bits_client_xact_id = RocketTile_1_io_uncached_0_acquire_bits_client_xact_id;
  assign uncore_io_tiles_uncached_0_acquire_bits_addr_beat = RocketTile_1_io_uncached_0_acquire_bits_addr_beat;
  assign uncore_io_tiles_uncached_0_acquire_bits_is_builtin_type = RocketTile_1_io_uncached_0_acquire_bits_is_builtin_type;
  assign uncore_io_tiles_uncached_0_acquire_bits_a_type = RocketTile_1_io_uncached_0_acquire_bits_a_type;
  assign uncore_io_tiles_uncached_0_acquire_bits_union = RocketTile_1_io_uncached_0_acquire_bits_union;
  assign uncore_io_tiles_uncached_0_acquire_bits_data = RocketTile_1_io_uncached_0_acquire_bits_data;
  assign uncore_io_tiles_uncached_0_grant_ready = RocketTile_1_io_uncached_0_grant_ready;
  assign uncore_io_mmio_axi_0_aw_ready = io_mmio_axi_0_aw_ready;
  assign uncore_io_mmio_axi_0_w_ready = io_mmio_axi_0_w_ready;
  assign uncore_io_mmio_axi_0_b_valid = io_mmio_axi_0_b_valid;
  assign uncore_io_mmio_axi_0_b_bits_resp = io_mmio_axi_0_b_bits_resp;
  assign uncore_io_mmio_axi_0_b_bits_id = io_mmio_axi_0_b_bits_id;
  assign uncore_io_mmio_axi_0_b_bits_user = io_mmio_axi_0_b_bits_user;
  assign uncore_io_mmio_axi_0_ar_ready = io_mmio_axi_0_ar_ready;
  assign uncore_io_mmio_axi_0_r_valid = io_mmio_axi_0_r_valid;
  assign uncore_io_mmio_axi_0_r_bits_resp = io_mmio_axi_0_r_bits_resp;
  assign uncore_io_mmio_axi_0_r_bits_data = io_mmio_axi_0_r_bits_data;
  assign uncore_io_mmio_axi_0_r_bits_last = io_mmio_axi_0_r_bits_last;
  assign uncore_io_mmio_axi_0_r_bits_id = io_mmio_axi_0_r_bits_id;
  assign uncore_io_mmio_axi_0_r_bits_user = io_mmio_axi_0_r_bits_user;
  assign uncore_io_interrupts_0 = io_interrupts_0;
  assign uncore_io_interrupts_1 = io_interrupts_1;
  assign uncore_io_interrupts_2 = io_interrupts_2;
  assign uncore_io_interrupts_3 = io_interrupts_3;
  assign uncore_io_interrupts_4 = io_interrupts_4;
  assign uncore_io_interrupts_5 = io_interrupts_5;
  assign uncore_io_interrupts_6 = io_interrupts_6;
  assign uncore_io_interrupts_7 = io_interrupts_7;
  assign uncore_io_interrupts_8 = io_interrupts_8;
  assign uncore_io_interrupts_9 = io_interrupts_9;
  assign uncore_io_interrupts_10 = io_interrupts_10;
  assign uncore_io_interrupts_11 = io_interrupts_11;
  assign uncore_io_interrupts_12 = io_interrupts_12;
  assign uncore_io_interrupts_13 = io_interrupts_13;
  assign uncore_io_interrupts_14 = io_interrupts_14;
  assign uncore_io_interrupts_15 = io_interrupts_15;
  assign uncore_io_interrupts_16 = io_interrupts_16;
  assign uncore_io_interrupts_17 = io_interrupts_17;
  assign uncore_io_interrupts_18 = io_interrupts_18;
  assign uncore_io_interrupts_19 = io_interrupts_19;
  assign uncore_io_interrupts_20 = io_interrupts_20;
  assign uncore_io_interrupts_21 = io_interrupts_21;
  assign uncore_io_interrupts_22 = io_interrupts_22;
  assign uncore_io_interrupts_23 = io_interrupts_23;
  assign uncore_io_interrupts_24 = io_interrupts_24;
  assign uncore_io_interrupts_25 = io_interrupts_25;
  assign uncore_io_interrupts_26 = io_interrupts_26;
  assign uncore_io_interrupts_27 = io_interrupts_27;
  assign uncore_io_interrupts_28 = io_interrupts_28;
  assign uncore_io_interrupts_29 = io_interrupts_29;
  assign uncore_io_interrupts_30 = io_interrupts_30;
  assign uncore_io_debugBus_req_valid = io_debug_req_valid;
  assign uncore_io_debugBus_req_bits_addr = io_debug_req_bits_addr;
  assign uncore_io_debugBus_req_bits_op = io_debug_req_bits_op;
  assign uncore_io_debugBus_req_bits_data = io_debug_req_bits_data;
  assign uncore_io_debugBus_resp_ready = io_debug_resp_ready;
endmodule
